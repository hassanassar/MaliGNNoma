`timescale 1 ps / 1 ps
`define XIL_TIMING

(* dont_touch = "true" *) 
(* NotValidForBitStream *)
module switch_elements
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  wire clk_i;
  wire [31:0]enable_i;
  (* DONT_TOUCH *) wire [31:0]info_s;
  wire rst_i;

  assign info_o[31:0] = info_s;
  (* DONT_TOUCH *) 
  (* NOISE_CIRC_AMOUNT = "7" *) 
  switch_elements_noise_source_wrapper \activity_blocks[0].switch 
       (.dummy_ext_signal(enable_i[1]),
        .dummy_output_o(info_s[0]),
        .loadseed_i(rst_i),
        .noise_enable_i(enable_i[0]),
        .randomize_active_instances(enable_i[2]),
        .sysclk(clk_i));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(info_s[31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(info_s[30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_s[21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_s[20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_s[19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_s[18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_s[17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_s[16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_s[15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_s[14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_s[13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_s[12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(info_s[29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_s[11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_s[10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_s[9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_s[8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_s[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_25
       (.I0(1'b0),
        .O(info_s[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_26
       (.I0(1'b0),
        .O(info_s[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_27
       (.I0(1'b0),
        .O(info_s[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_28
       (.I0(1'b0),
        .O(info_s[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_29
       (.I0(1'b0),
        .O(info_s[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(info_s[28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_30
       (.I0(1'b0),
        .O(info_s[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(info_s[27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(info_s[26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(info_s[25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(info_s[24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(info_s[23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_s[22]));
endmodule

(* NOISE_CIRC_AMOUNT = "7" *) (* ORIG_REF_NAME = "noise_source_wrapper" *) (* dont_touch = "true" *) 
module switch_elements_noise_source_wrapper
   (sysclk,
    loadseed_i,
    noise_enable_i,
    dummy_ext_signal,
    dummy_output_o,
    randomize_active_instances);
  input sysclk;
  input loadseed_i;
  input noise_enable_i;
  input dummy_ext_signal;
  output dummy_output_o;
  input randomize_active_instances;

  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[0] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[1] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[2] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[3] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[4] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[5] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [30:0]\bench_v[6] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[0] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[1] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[2] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[3] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[4] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[5] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout[6] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[0] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[1] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[2] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[3] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[4] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[5] ;
  (* DONT_TOUCH *) (* MARK_DEBUG *) (* RTL_KEEP = "true" *) 
  (* S *) wire [120:0]\bench_vout_reg[6] ;
  wire clear;
  wire dummy_output_o;
  wire \en_counter[8]_i_3_n_0 ;
  wire \en_counter[8]_i_4_n_0 ;
  wire [0:0]en_counter_reg;
  wire [8:1]en_counter_reg__0;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) wire loadseed_s;
  wire n_noise_enable_s;
  (* RTL_KEEP = "true" *) wire noise_enable_s;
  wire [8:0]plusOp;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[0] ;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[1] ;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[2] ;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[3] ;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[4] ;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[5] ;
  (* MARK_DEBUG *) (* RTL_KEEP = "true" *) (* S *) wire [31:0]\random_data_s[6] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[0] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[1] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[2] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[3] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[4] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[5] ;
  (* RTL_KEEP = "true" *) (* S *) wire [31:0]\seed_s[6] ;
  wire sysclk;

  assign loadseed_s = loadseed_i;
  assign noise_enable_s = noise_enable_i;
  assign \seed_s[6] [0] = dummy_ext_signal;
  LUT3 #(
    .INIT(8'hB8)) 
    dummy_output_o_INST_0
       (.I0(\bench_vout_reg[1] [1]),
        .I1(en_counter_reg),
        .I2(\bench_vout_reg[0] [0]),
        .O(dummy_output_o));
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \en_counter[0]_i_1 
       (.I0(en_counter_reg),
        .O(plusOp[0]));
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \en_counter[1]_i_1 
       (.I0(en_counter_reg),
        .I1(en_counter_reg__0[1]),
        .O(plusOp[1]));
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \en_counter[2]_i_1 
       (.I0(en_counter_reg),
        .I1(en_counter_reg__0[1]),
        .I2(en_counter_reg__0[2]),
        .O(plusOp[2]));
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \en_counter[3]_i_1 
       (.I0(en_counter_reg__0[1]),
        .I1(en_counter_reg),
        .I2(en_counter_reg__0[2]),
        .I3(en_counter_reg__0[3]),
        .O(plusOp[3]));
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \en_counter[4]_i_1 
       (.I0(en_counter_reg__0[2]),
        .I1(en_counter_reg),
        .I2(en_counter_reg__0[1]),
        .I3(en_counter_reg__0[3]),
        .I4(en_counter_reg__0[4]),
        .O(plusOp[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \en_counter[5]_i_1 
       (.I0(en_counter_reg__0[3]),
        .I1(en_counter_reg__0[1]),
        .I2(en_counter_reg),
        .I3(en_counter_reg__0[2]),
        .I4(en_counter_reg__0[4]),
        .I5(en_counter_reg__0[5]),
        .O(plusOp[5]));
  LUT2 #(
    .INIT(4'h6)) 
    \en_counter[6]_i_1 
       (.I0(\en_counter[8]_i_4_n_0 ),
        .I1(en_counter_reg__0[6]),
        .O(plusOp[6]));
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \en_counter[7]_i_1 
       (.I0(\en_counter[8]_i_4_n_0 ),
        .I1(en_counter_reg__0[6]),
        .I2(en_counter_reg__0[7]),
        .O(plusOp[7]));
  LUT5 #(
    .INIT(32'hAAA8AAAA)) 
    \en_counter[8]_i_1 
       (.I0(en_counter_reg__0[8]),
        .I1(en_counter_reg__0[5]),
        .I2(en_counter_reg__0[7]),
        .I3(en_counter_reg__0[6]),
        .I4(\en_counter[8]_i_3_n_0 ),
        .O(clear));
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \en_counter[8]_i_2 
       (.I0(en_counter_reg__0[6]),
        .I1(\en_counter[8]_i_4_n_0 ),
        .I2(en_counter_reg__0[7]),
        .I3(en_counter_reg__0[8]),
        .O(plusOp[8]));
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT5 #(
    .INIT(32'h0155FFFF)) 
    \en_counter[8]_i_3 
       (.I0(en_counter_reg__0[3]),
        .I1(en_counter_reg),
        .I2(en_counter_reg__0[1]),
        .I3(en_counter_reg__0[2]),
        .I4(en_counter_reg__0[4]),
        .O(\en_counter[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \en_counter[8]_i_4 
       (.I0(en_counter_reg__0[5]),
        .I1(en_counter_reg__0[3]),
        .I2(en_counter_reg__0[1]),
        .I3(en_counter_reg),
        .I4(en_counter_reg__0[2]),
        .I5(en_counter_reg__0[4]),
        .O(\en_counter[8]_i_4_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[0]),
        .Q(en_counter_reg),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[1]),
        .Q(en_counter_reg__0[1]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[2]),
        .Q(en_counter_reg__0[2]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[3]),
        .Q(en_counter_reg__0[3]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[4]),
        .Q(en_counter_reg__0[4]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[5]),
        .Q(en_counter_reg__0[5]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[6]),
        .Q(en_counter_reg__0[6]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[7]),
        .Q(en_counter_reg__0[7]),
        .R(clear));
  FDRE #(
    .INIT(1'b0)) 
    \en_counter_reg[8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(plusOp[8]),
        .Q(en_counter_reg__0[8]),
        .R(clear));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(\seed_s[1] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(\seed_s[1] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(\seed_s[1] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_100
       (.I0(1'b0),
        .O(\seed_s[3] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_101
       (.I0(1'b0),
        .O(\seed_s[3] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_102
       (.I0(1'b0),
        .O(\seed_s[3] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_103
       (.I0(1'b0),
        .O(\seed_s[3] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_104
       (.I0(1'b0),
        .O(\seed_s[3] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_105
       (.I0(1'b1),
        .O(\seed_s[3] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_106
       (.I0(1'b0),
        .O(\seed_s[3] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_107
       (.I0(1'b0),
        .O(\seed_s[3] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_108
       (.I0(1'b0),
        .O(\seed_s[3] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_109
       (.I0(1'b0),
        .O(\seed_s[3] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(\seed_s[1] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_110
       (.I0(1'b0),
        .O(\seed_s[3] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_111
       (.I0(1'b0),
        .O(\seed_s[3] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_112
       (.I0(1'b0),
        .O(\seed_s[3] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_113
       (.I0(1'b0),
        .O(\seed_s[3] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_114
       (.I0(1'b0),
        .O(\seed_s[3] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_115
       (.I0(1'b0),
        .O(\seed_s[3] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_116
       (.I0(1'b0),
        .O(\seed_s[3] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_117
       (.I0(1'b0),
        .O(\seed_s[3] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_118
       (.I0(1'b0),
        .O(\seed_s[3] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_119
       (.I0(1'b0),
        .O(\seed_s[3] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(\seed_s[1] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_120
       (.I0(1'b0),
        .O(\seed_s[3] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_121
       (.I0(1'b1),
        .O(\seed_s[3] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_122
       (.I0(1'b0),
        .O(\seed_s[3] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_123
       (.I0(1'b0),
        .O(\seed_s[3] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_124
       (.I0(1'b0),
        .O(\seed_s[4] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_125
       (.I0(1'b0),
        .O(\seed_s[4] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_126
       (.I0(1'b0),
        .O(\seed_s[4] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_127
       (.I0(1'b0),
        .O(\seed_s[4] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_128
       (.I0(1'b0),
        .O(\seed_s[4] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_129
       (.I0(1'b0),
        .O(\seed_s[4] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b1),
        .O(\seed_s[1] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_130
       (.I0(1'b0),
        .O(\seed_s[4] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_131
       (.I0(1'b0),
        .O(\seed_s[4] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_132
       (.I0(1'b0),
        .O(\seed_s[4] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_133
       (.I0(1'b0),
        .O(\seed_s[4] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_134
       (.I0(1'b0),
        .O(\seed_s[4] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_135
       (.I0(1'b0),
        .O(\seed_s[4] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_136
       (.I0(1'b1),
        .O(\seed_s[4] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_137
       (.I0(1'b0),
        .O(\seed_s[4] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_138
       (.I0(1'b1),
        .O(\seed_s[4] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_139
       (.I0(1'b0),
        .O(\seed_s[4] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(\seed_s[1] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_140
       (.I0(1'b0),
        .O(\seed_s[4] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_141
       (.I0(1'b0),
        .O(\seed_s[4] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_142
       (.I0(1'b0),
        .O(\seed_s[4] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_143
       (.I0(1'b0),
        .O(\seed_s[4] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_144
       (.I0(1'b0),
        .O(\seed_s[4] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_145
       (.I0(1'b0),
        .O(\seed_s[4] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_146
       (.I0(1'b0),
        .O(\seed_s[4] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_147
       (.I0(1'b0),
        .O(\seed_s[4] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_148
       (.I0(1'b0),
        .O(\seed_s[4] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_149
       (.I0(1'b0),
        .O(\seed_s[4] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(\seed_s[1] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_150
       (.I0(1'b0),
        .O(\seed_s[4] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_151
       (.I0(1'b0),
        .O(\seed_s[4] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_152
       (.I0(1'b1),
        .O(\seed_s[4] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_153
       (.I0(1'b0),
        .O(\seed_s[4] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_154
       (.I0(1'b1),
        .O(\seed_s[4] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_155
       (.I0(1'b0),
        .O(\seed_s[5] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_156
       (.I0(1'b0),
        .O(\seed_s[5] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_157
       (.I0(1'b0),
        .O(\seed_s[5] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_158
       (.I0(1'b0),
        .O(\seed_s[5] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_159
       (.I0(1'b0),
        .O(\seed_s[5] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(\seed_s[1] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_160
       (.I0(1'b0),
        .O(\seed_s[5] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_161
       (.I0(1'b0),
        .O(\seed_s[5] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_162
       (.I0(1'b0),
        .O(\seed_s[5] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_163
       (.I0(1'b0),
        .O(\seed_s[5] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_164
       (.I0(1'b0),
        .O(\seed_s[5] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_165
       (.I0(1'b0),
        .O(\seed_s[5] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_166
       (.I0(1'b0),
        .O(\seed_s[5] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_167
       (.I0(1'b1),
        .O(\seed_s[5] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_168
       (.I0(1'b1),
        .O(\seed_s[5] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_169
       (.I0(1'b0),
        .O(\seed_s[5] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(\seed_s[1] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_170
       (.I0(1'b0),
        .O(\seed_s[5] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_171
       (.I0(1'b0),
        .O(\seed_s[5] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_172
       (.I0(1'b0),
        .O(\seed_s[5] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_173
       (.I0(1'b0),
        .O(\seed_s[5] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_174
       (.I0(1'b0),
        .O(\seed_s[5] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_175
       (.I0(1'b0),
        .O(\seed_s[5] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_176
       (.I0(1'b0),
        .O(\seed_s[5] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_177
       (.I0(1'b0),
        .O(\seed_s[5] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_178
       (.I0(1'b0),
        .O(\seed_s[5] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_179
       (.I0(1'b0),
        .O(\seed_s[5] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(\seed_s[1] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_180
       (.I0(1'b0),
        .O(\seed_s[5] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_181
       (.I0(1'b0),
        .O(\seed_s[5] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_182
       (.I0(1'b0),
        .O(\seed_s[5] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_183
       (.I0(1'b1),
        .O(\seed_s[5] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_184
       (.I0(1'b1),
        .O(\seed_s[5] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_185
       (.I0(1'b0),
        .O(\seed_s[5] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_186
       (.I0(1'b0),
        .O(\seed_s[6] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_187
       (.I0(1'b0),
        .O(\seed_s[6] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_188
       (.I0(1'b0),
        .O(\seed_s[6] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_189
       (.I0(1'b0),
        .O(\seed_s[6] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(\seed_s[1] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_190
       (.I0(1'b0),
        .O(\seed_s[6] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_191
       (.I0(1'b0),
        .O(\seed_s[6] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_192
       (.I0(1'b0),
        .O(\seed_s[6] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_193
       (.I0(1'b0),
        .O(\seed_s[6] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_194
       (.I0(1'b0),
        .O(\seed_s[6] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_195
       (.I0(1'b0),
        .O(\seed_s[6] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_196
       (.I0(1'b0),
        .O(\seed_s[6] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_197
       (.I0(1'b0),
        .O(\seed_s[6] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_198
       (.I0(1'b1),
        .O(\seed_s[6] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_199
       (.I0(1'b1),
        .O(\seed_s[6] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(\seed_s[1] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(\seed_s[1] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_200
       (.I0(1'b1),
        .O(\seed_s[6] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_201
       (.I0(1'b0),
        .O(\seed_s[6] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_202
       (.I0(1'b0),
        .O(\seed_s[6] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_203
       (.I0(1'b0),
        .O(\seed_s[6] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_204
       (.I0(1'b0),
        .O(\seed_s[6] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_205
       (.I0(1'b0),
        .O(\seed_s[6] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_206
       (.I0(1'b0),
        .O(\seed_s[6] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_207
       (.I0(1'b0),
        .O(\seed_s[6] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_208
       (.I0(1'b0),
        .O(\seed_s[6] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_209
       (.I0(1'b0),
        .O(\seed_s[6] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(\seed_s[1] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_210
       (.I0(1'b0),
        .O(\seed_s[6] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_211
       (.I0(1'b0),
        .O(\seed_s[6] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_212
       (.I0(1'b0),
        .O(\seed_s[6] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_213
       (.I0(1'b0),
        .O(\seed_s[6] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_214
       (.I0(1'b1),
        .O(\seed_s[6] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_215
       (.I0(1'b1),
        .O(\seed_s[6] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_216
       (.I0(1'b1),
        .O(\seed_s[6] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(\seed_s[1] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(\seed_s[1] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(\seed_s[1] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_25
       (.I0(1'b0),
        .O(\seed_s[1] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_26
       (.I0(1'b0),
        .O(\seed_s[1] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_27
       (.I0(1'b0),
        .O(\seed_s[1] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_28
       (.I0(1'b0),
        .O(\seed_s[1] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_29
       (.I0(1'b1),
        .O(\seed_s[1] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(\seed_s[1] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_30
       (.I0(1'b0),
        .O(\seed_s[1] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_31
       (.I0(1'b0),
        .O(\seed_s[0] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_32
       (.I0(1'b0),
        .O(\seed_s[0] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_33
       (.I0(1'b0),
        .O(\seed_s[0] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_34
       (.I0(1'b0),
        .O(\seed_s[0] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_35
       (.I0(1'b0),
        .O(\seed_s[0] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_36
       (.I0(1'b0),
        .O(\seed_s[0] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_37
       (.I0(1'b0),
        .O(\seed_s[0] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_38
       (.I0(1'b0),
        .O(\seed_s[0] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_39
       (.I0(1'b0),
        .O(\seed_s[0] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(\seed_s[1] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_40
       (.I0(1'b0),
        .O(\seed_s[0] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_41
       (.I0(1'b0),
        .O(\seed_s[0] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_42
       (.I0(1'b0),
        .O(\seed_s[0] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_43
       (.I0(1'b0),
        .O(\seed_s[0] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_44
       (.I0(1'b0),
        .O(\seed_s[0] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_45
       (.I0(1'b1),
        .O(\seed_s[0] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_46
       (.I0(1'b0),
        .O(\seed_s[0] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_47
       (.I0(1'b0),
        .O(\seed_s[0] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_48
       (.I0(1'b0),
        .O(\seed_s[0] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_49
       (.I0(1'b0),
        .O(\seed_s[0] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(\seed_s[1] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_50
       (.I0(1'b0),
        .O(\seed_s[0] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_51
       (.I0(1'b0),
        .O(\seed_s[0] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_52
       (.I0(1'b0),
        .O(\seed_s[0] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_53
       (.I0(1'b0),
        .O(\seed_s[0] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_54
       (.I0(1'b0),
        .O(\seed_s[0] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_55
       (.I0(1'b0),
        .O(\seed_s[0] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_56
       (.I0(1'b0),
        .O(\seed_s[0] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_57
       (.I0(1'b0),
        .O(\seed_s[0] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_58
       (.I0(1'b0),
        .O(\seed_s[0] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_59
       (.I0(1'b0),
        .O(\seed_s[0] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(\seed_s[1] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_60
       (.I0(1'b0),
        .O(\seed_s[0] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_61
       (.I0(1'b1),
        .O(\seed_s[0] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_62
       (.I0(1'b0),
        .O(\seed_s[2] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_63
       (.I0(1'b0),
        .O(\seed_s[2] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_64
       (.I0(1'b0),
        .O(\seed_s[2] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_65
       (.I0(1'b0),
        .O(\seed_s[2] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_66
       (.I0(1'b0),
        .O(\seed_s[2] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_67
       (.I0(1'b0),
        .O(\seed_s[2] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_68
       (.I0(1'b0),
        .O(\seed_s[2] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    i_69
       (.I0(1'b0),
        .O(\seed_s[2] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(\seed_s[1] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    i_70
       (.I0(1'b0),
        .O(\seed_s[2] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_71
       (.I0(1'b0),
        .O(\seed_s[2] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_72
       (.I0(1'b0),
        .O(\seed_s[2] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    i_73
       (.I0(1'b0),
        .O(\seed_s[2] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    i_74
       (.I0(1'b0),
        .O(\seed_s[2] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    i_75
       (.I0(1'b1),
        .O(\seed_s[2] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_76
       (.I0(1'b1),
        .O(\seed_s[2] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    i_77
       (.I0(1'b0),
        .O(\seed_s[2] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    i_78
       (.I0(1'b0),
        .O(\seed_s[2] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_79
       (.I0(1'b0),
        .O(\seed_s[2] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(\seed_s[1] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    i_80
       (.I0(1'b0),
        .O(\seed_s[2] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_81
       (.I0(1'b0),
        .O(\seed_s[2] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_82
       (.I0(1'b0),
        .O(\seed_s[2] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_83
       (.I0(1'b0),
        .O(\seed_s[2] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_84
       (.I0(1'b0),
        .O(\seed_s[2] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_85
       (.I0(1'b0),
        .O(\seed_s[2] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_86
       (.I0(1'b0),
        .O(\seed_s[2] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_87
       (.I0(1'b0),
        .O(\seed_s[2] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_88
       (.I0(1'b0),
        .O(\seed_s[2] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_89
       (.I0(1'b0),
        .O(\seed_s[2] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(\seed_s[1] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    i_90
       (.I0(1'b0),
        .O(\seed_s[2] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_91
       (.I0(1'b1),
        .O(\seed_s[2] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_92
       (.I0(1'b1),
        .O(\seed_s[2] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_93
       (.I0(1'b0),
        .O(\seed_s[3] [31]));
  LUT1 #(
    .INIT(2'h2)) 
    i_94
       (.I0(1'b0),
        .O(\seed_s[3] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    i_95
       (.I0(1'b0),
        .O(\seed_s[3] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    i_96
       (.I0(1'b0),
        .O(\seed_s[3] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    i_97
       (.I0(1'b0),
        .O(\seed_s[3] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    i_98
       (.I0(1'b0),
        .O(\seed_s[3] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    i_99
       (.I0(1'b0),
        .O(\seed_s[3] [25]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [0]),
        .Q(\bench_vout_reg[0] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [100]),
        .Q(\bench_vout_reg[0] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [101]),
        .Q(\bench_vout_reg[0] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [102]),
        .Q(\bench_vout_reg[0] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [103]),
        .Q(\bench_vout_reg[0] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [104]),
        .Q(\bench_vout_reg[0] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [105]),
        .Q(\bench_vout_reg[0] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [106]),
        .Q(\bench_vout_reg[0] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [107]),
        .Q(\bench_vout_reg[0] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [108]),
        .Q(\bench_vout_reg[0] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [109]),
        .Q(\bench_vout_reg[0] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [10]),
        .Q(\bench_vout_reg[0] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [110]),
        .Q(\bench_vout_reg[0] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [111]),
        .Q(\bench_vout_reg[0] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [112]),
        .Q(\bench_vout_reg[0] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [113]),
        .Q(\bench_vout_reg[0] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [114]),
        .Q(\bench_vout_reg[0] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [115]),
        .Q(\bench_vout_reg[0] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [116]),
        .Q(\bench_vout_reg[0] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [117]),
        .Q(\bench_vout_reg[0] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [118]),
        .Q(\bench_vout_reg[0] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [119]),
        .Q(\bench_vout_reg[0] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [11]),
        .Q(\bench_vout_reg[0] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [120]),
        .Q(\bench_vout_reg[0] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [12]),
        .Q(\bench_vout_reg[0] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [13]),
        .Q(\bench_vout_reg[0] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [14]),
        .Q(\bench_vout_reg[0] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [15]),
        .Q(\bench_vout_reg[0] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [16]),
        .Q(\bench_vout_reg[0] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [17]),
        .Q(\bench_vout_reg[0] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [18]),
        .Q(\bench_vout_reg[0] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [19]),
        .Q(\bench_vout_reg[0] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [1]),
        .Q(\bench_vout_reg[0] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [20]),
        .Q(\bench_vout_reg[0] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [21]),
        .Q(\bench_vout_reg[0] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [22]),
        .Q(\bench_vout_reg[0] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [23]),
        .Q(\bench_vout_reg[0] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [24]),
        .Q(\bench_vout_reg[0] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [25]),
        .Q(\bench_vout_reg[0] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [26]),
        .Q(\bench_vout_reg[0] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [27]),
        .Q(\bench_vout_reg[0] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [28]),
        .Q(\bench_vout_reg[0] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [29]),
        .Q(\bench_vout_reg[0] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [2]),
        .Q(\bench_vout_reg[0] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [30]),
        .Q(\bench_vout_reg[0] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [31]),
        .Q(\bench_vout_reg[0] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [32]),
        .Q(\bench_vout_reg[0] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [33]),
        .Q(\bench_vout_reg[0] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [34]),
        .Q(\bench_vout_reg[0] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [35]),
        .Q(\bench_vout_reg[0] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [36]),
        .Q(\bench_vout_reg[0] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [37]),
        .Q(\bench_vout_reg[0] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [38]),
        .Q(\bench_vout_reg[0] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [39]),
        .Q(\bench_vout_reg[0] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [3]),
        .Q(\bench_vout_reg[0] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [40]),
        .Q(\bench_vout_reg[0] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [41]),
        .Q(\bench_vout_reg[0] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [42]),
        .Q(\bench_vout_reg[0] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [43]),
        .Q(\bench_vout_reg[0] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [44]),
        .Q(\bench_vout_reg[0] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [45]),
        .Q(\bench_vout_reg[0] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [46]),
        .Q(\bench_vout_reg[0] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [47]),
        .Q(\bench_vout_reg[0] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [48]),
        .Q(\bench_vout_reg[0] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [49]),
        .Q(\bench_vout_reg[0] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [4]),
        .Q(\bench_vout_reg[0] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [50]),
        .Q(\bench_vout_reg[0] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [51]),
        .Q(\bench_vout_reg[0] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [52]),
        .Q(\bench_vout_reg[0] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [53]),
        .Q(\bench_vout_reg[0] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [54]),
        .Q(\bench_vout_reg[0] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [55]),
        .Q(\bench_vout_reg[0] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [56]),
        .Q(\bench_vout_reg[0] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [57]),
        .Q(\bench_vout_reg[0] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [58]),
        .Q(\bench_vout_reg[0] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [59]),
        .Q(\bench_vout_reg[0] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [5]),
        .Q(\bench_vout_reg[0] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [60]),
        .Q(\bench_vout_reg[0] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [61]),
        .Q(\bench_vout_reg[0] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [62]),
        .Q(\bench_vout_reg[0] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [63]),
        .Q(\bench_vout_reg[0] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [64]),
        .Q(\bench_vout_reg[0] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [65]),
        .Q(\bench_vout_reg[0] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [66]),
        .Q(\bench_vout_reg[0] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [67]),
        .Q(\bench_vout_reg[0] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [68]),
        .Q(\bench_vout_reg[0] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [69]),
        .Q(\bench_vout_reg[0] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [6]),
        .Q(\bench_vout_reg[0] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [70]),
        .Q(\bench_vout_reg[0] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [71]),
        .Q(\bench_vout_reg[0] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [72]),
        .Q(\bench_vout_reg[0] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [73]),
        .Q(\bench_vout_reg[0] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [74]),
        .Q(\bench_vout_reg[0] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [75]),
        .Q(\bench_vout_reg[0] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [76]),
        .Q(\bench_vout_reg[0] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [77]),
        .Q(\bench_vout_reg[0] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [78]),
        .Q(\bench_vout_reg[0] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [79]),
        .Q(\bench_vout_reg[0] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [7]),
        .Q(\bench_vout_reg[0] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [80]),
        .Q(\bench_vout_reg[0] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [81]),
        .Q(\bench_vout_reg[0] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [82]),
        .Q(\bench_vout_reg[0] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [83]),
        .Q(\bench_vout_reg[0] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [84]),
        .Q(\bench_vout_reg[0] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [85]),
        .Q(\bench_vout_reg[0] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [86]),
        .Q(\bench_vout_reg[0] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [87]),
        .Q(\bench_vout_reg[0] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [88]),
        .Q(\bench_vout_reg[0] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [89]),
        .Q(\bench_vout_reg[0] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [8]),
        .Q(\bench_vout_reg[0] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [90]),
        .Q(\bench_vout_reg[0] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [91]),
        .Q(\bench_vout_reg[0] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [92]),
        .Q(\bench_vout_reg[0] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [93]),
        .Q(\bench_vout_reg[0] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [94]),
        .Q(\bench_vout_reg[0] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [95]),
        .Q(\bench_vout_reg[0] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [96]),
        .Q(\bench_vout_reg[0] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [97]),
        .Q(\bench_vout_reg[0] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [98]),
        .Q(\bench_vout_reg[0] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [99]),
        .Q(\bench_vout_reg[0] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[0].bench_vout_reg_reg[0][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[0] [9]),
        .Q(\bench_vout_reg[0] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng__1 \noise_circ_replica[0].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[0] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[0] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench__1 \noise_circ_replica[0].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[0] [24]),
        .g1006(\bench_vout[0] [7]),
        .g1008(\bench_v[0] [25]),
        .g1015(\bench_vout[0] [8]),
        .g1016(\bench_v[0] [26]),
        .g1017(\bench_vout[0] [9]),
        .g1080(\bench_v[0] [27]),
        .g1234(\bench_v[0] [28]),
        .g1246(\bench_vout[0] [10]),
        .g1553(\bench_v[0] [29]),
        .g1554(\bench_v[0] [30]),
        .g1724(\bench_vout[0] [11]),
        .g1783(\bench_vout[0] [12]),
        .g1798(\bench_vout[0] [13]),
        .g1804(\bench_vout[0] [14]),
        .g1810(\bench_vout[0] [15]),
        .g1817(\bench_vout[0] [16]),
        .g1824(\bench_vout[0] [17]),
        .g1829(\bench_vout[0] [18]),
        .g1870(\bench_vout[0] [19]),
        .g1871(\bench_vout[0] [20]),
        .g1894(\bench_vout[0] [21]),
        .g1911(\bench_vout[0] [22]),
        .g1944(\bench_vout[0] [23]),
        .g206(\bench_vout[0] [0]),
        .g2662(\bench_vout[0] [24]),
        .g2844(\bench_vout[0] [25]),
        .g2888(\bench_vout[0] [26]),
        .g291(\bench_vout[0] [1]),
        .g3077(\bench_vout[0] [27]),
        .g3096(\bench_vout[0] [28]),
        .g3130(\bench_vout[0] [29]),
        .g3159(\bench_vout[0] [30]),
        .g3191(\bench_vout[0] [31]),
        .g372(\bench_vout[0] [2]),
        .g3829(\bench_vout[0] [32]),
        .g3859(\bench_vout[0] [33]),
        .g3860(\bench_vout[0] [34]),
        .g4267(\bench_vout[0] [35]),
        .g43(\bench_v[0] [0]),
        .g4316(\bench_vout[0] [36]),
        .g4370(\bench_vout[0] [37]),
        .g4371(\bench_vout[0] [38]),
        .g4372(\bench_vout[0] [39]),
        .g4373(\bench_vout[0] [40]),
        .g453(\bench_vout[0] [3]),
        .g4655(\bench_vout[0] [41]),
        .g4657(\bench_vout[0] [42]),
        .g4660(\bench_vout[0] [43]),
        .g4661(\bench_vout[0] [44]),
        .g4663(\bench_vout[0] [45]),
        .g4664(\bench_vout[0] [46]),
        .g49(\bench_v[0] [1]),
        .g5143(\bench_vout[0] [47]),
        .g5164(\bench_vout[0] [48]),
        .g534(\bench_vout[0] [4]),
        .g5571(\bench_vout[0] [49]),
        .g5669(\bench_vout[0] [50]),
        .g5678(\bench_vout[0] [51]),
        .g5682(\bench_vout[0] [52]),
        .g5684(\bench_vout[0] [53]),
        .g5687(\bench_vout[0] [54]),
        .g5729(\bench_vout[0] [55]),
        .g594(\bench_vout[0] [5]),
        .g6207(\bench_vout[0] [56]),
        .g6212(\bench_vout[0] [57]),
        .g6223(\bench_vout[0] [58]),
        .g6236(\bench_vout[0] [59]),
        .g6269(\bench_vout[0] [60]),
        .g633(\bench_v[0] [2]),
        .g634(\bench_v[0] [3]),
        .g635(\bench_v[0] [4]),
        .g6425(\bench_vout[0] [61]),
        .g645(\bench_v[0] [5]),
        .g647(\bench_v[0] [6]),
        .g648(\bench_v[0] [7]),
        .g6648(\bench_vout[0] [62]),
        .g6653(\bench_vout[0] [63]),
        .g6675(\bench_vout[0] [64]),
        .g6849(\bench_vout[0] [65]),
        .g6850(\bench_vout[0] [66]),
        .g6895(\bench_vout[0] [67]),
        .g690(\bench_v[0] [8]),
        .g6909(\bench_vout[0] [68]),
        .g694(\bench_v[0] [9]),
        .g698(\bench_v[0] [10]),
        .g702(\bench_v[0] [11]),
        .g7048(\bench_vout[0] [69]),
        .g7063(\bench_vout[0] [70]),
        .g7103(\bench_vout[0] [71]),
        .g722(\bench_v[0] [12]),
        .g723(\bench_v[0] [13]),
        .g7283(\bench_vout[0] [72]),
        .g7284(\bench_vout[0] [73]),
        .g7285(\bench_vout[0] [74]),
        .g7286(\bench_vout[0] [75]),
        .g7287(\bench_vout[0] [76]),
        .g7288(\bench_vout[0] [77]),
        .g7289(\bench_vout[0] [78]),
        .g7290(\bench_vout[0] [79]),
        .g7291(\bench_vout[0] [80]),
        .g7292(\bench_vout[0] [81]),
        .g7293(\bench_vout[0] [82]),
        .g7294(\bench_vout[0] [83]),
        .g7295(\bench_vout[0] [84]),
        .g7298(\bench_vout[0] [85]),
        .g7423(\bench_vout[0] [86]),
        .g7424(\bench_vout[0] [87]),
        .g7425(\bench_vout[0] [88]),
        .g7474(\bench_vout[0] [89]),
        .g7504(\bench_vout[0] [90]),
        .g7505(\bench_vout[0] [91]),
        .g7506(\bench_vout[0] [92]),
        .g7507(\bench_vout[0] [93]),
        .g7508(\bench_vout[0] [94]),
        .g751(\bench_v[0] [14]),
        .g7514(\bench_vout[0] [95]),
        .g752(\bench_v[0] [15]),
        .g753(\bench_v[0] [16]),
        .g754(\bench_v[0] [17]),
        .g755(\bench_v[0] [18]),
        .g756(\bench_v[0] [19]),
        .g757(\bench_v[0] [20]),
        .g7729(\bench_vout[0] [96]),
        .g7730(\bench_vout[0] [97]),
        .g7731(\bench_vout[0] [98]),
        .g7732(\bench_vout[0] [99]),
        .g781(\bench_v[0] [21]),
        .g785(\bench_vout[0] [6]),
        .g8216(\bench_vout[0] [100]),
        .g8217(\bench_vout[0] [101]),
        .g8218(\bench_vout[0] [102]),
        .g8219(\bench_vout[0] [103]),
        .g8234(\bench_vout[0] [104]),
        .g8661(\bench_vout[0] [105]),
        .g8663(\bench_vout[0] [106]),
        .g8872(\bench_vout[0] [107]),
        .g8958(\bench_vout[0] [108]),
        .g9128(\bench_vout[0] [109]),
        .g9132(\bench_vout[0] [110]),
        .g9204(\bench_vout[0] [111]),
        .g9280(\bench_vout[0] [112]),
        .g9297(\bench_vout[0] [113]),
        .g9299(\bench_vout[0] [114]),
        .g9305(\bench_vout[0] [115]),
        .g9308(\bench_vout[0] [116]),
        .g9310(\bench_vout[0] [117]),
        .g9312(\bench_vout[0] [118]),
        .g9314(\bench_vout[0] [119]),
        .g9378(\bench_vout[0] [120]),
        .g941(\bench_v[0] [22]),
        .g962(\bench_v[0] [23]));
  LUT1 #(
    .INIT(2'h1)) 
    \noise_circ_replica[0].s13207_bench_inst_i_1 
       (.I0(noise_enable_s),
        .O(n_noise_enable_s));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [0]),
        .Q(\bench_vout_reg[1] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [100]),
        .Q(\bench_vout_reg[1] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [101]),
        .Q(\bench_vout_reg[1] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [102]),
        .Q(\bench_vout_reg[1] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [103]),
        .Q(\bench_vout_reg[1] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [104]),
        .Q(\bench_vout_reg[1] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [105]),
        .Q(\bench_vout_reg[1] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [106]),
        .Q(\bench_vout_reg[1] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [107]),
        .Q(\bench_vout_reg[1] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [108]),
        .Q(\bench_vout_reg[1] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [109]),
        .Q(\bench_vout_reg[1] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [10]),
        .Q(\bench_vout_reg[1] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [110]),
        .Q(\bench_vout_reg[1] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [111]),
        .Q(\bench_vout_reg[1] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [112]),
        .Q(\bench_vout_reg[1] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [113]),
        .Q(\bench_vout_reg[1] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [114]),
        .Q(\bench_vout_reg[1] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [115]),
        .Q(\bench_vout_reg[1] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [116]),
        .Q(\bench_vout_reg[1] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [117]),
        .Q(\bench_vout_reg[1] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [118]),
        .Q(\bench_vout_reg[1] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [119]),
        .Q(\bench_vout_reg[1] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [11]),
        .Q(\bench_vout_reg[1] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [120]),
        .Q(\bench_vout_reg[1] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [12]),
        .Q(\bench_vout_reg[1] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [13]),
        .Q(\bench_vout_reg[1] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [14]),
        .Q(\bench_vout_reg[1] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [15]),
        .Q(\bench_vout_reg[1] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [16]),
        .Q(\bench_vout_reg[1] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [17]),
        .Q(\bench_vout_reg[1] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [18]),
        .Q(\bench_vout_reg[1] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [19]),
        .Q(\bench_vout_reg[1] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [1]),
        .Q(\bench_vout_reg[1] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [20]),
        .Q(\bench_vout_reg[1] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [21]),
        .Q(\bench_vout_reg[1] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [22]),
        .Q(\bench_vout_reg[1] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [23]),
        .Q(\bench_vout_reg[1] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [24]),
        .Q(\bench_vout_reg[1] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [25]),
        .Q(\bench_vout_reg[1] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [26]),
        .Q(\bench_vout_reg[1] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [27]),
        .Q(\bench_vout_reg[1] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [28]),
        .Q(\bench_vout_reg[1] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [29]),
        .Q(\bench_vout_reg[1] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [2]),
        .Q(\bench_vout_reg[1] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [30]),
        .Q(\bench_vout_reg[1] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [31]),
        .Q(\bench_vout_reg[1] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [32]),
        .Q(\bench_vout_reg[1] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [33]),
        .Q(\bench_vout_reg[1] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [34]),
        .Q(\bench_vout_reg[1] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [35]),
        .Q(\bench_vout_reg[1] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [36]),
        .Q(\bench_vout_reg[1] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [37]),
        .Q(\bench_vout_reg[1] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [38]),
        .Q(\bench_vout_reg[1] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [39]),
        .Q(\bench_vout_reg[1] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [3]),
        .Q(\bench_vout_reg[1] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [40]),
        .Q(\bench_vout_reg[1] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [41]),
        .Q(\bench_vout_reg[1] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [42]),
        .Q(\bench_vout_reg[1] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [43]),
        .Q(\bench_vout_reg[1] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [44]),
        .Q(\bench_vout_reg[1] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [45]),
        .Q(\bench_vout_reg[1] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [46]),
        .Q(\bench_vout_reg[1] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [47]),
        .Q(\bench_vout_reg[1] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [48]),
        .Q(\bench_vout_reg[1] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [49]),
        .Q(\bench_vout_reg[1] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [4]),
        .Q(\bench_vout_reg[1] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [50]),
        .Q(\bench_vout_reg[1] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [51]),
        .Q(\bench_vout_reg[1] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [52]),
        .Q(\bench_vout_reg[1] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [53]),
        .Q(\bench_vout_reg[1] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [54]),
        .Q(\bench_vout_reg[1] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [55]),
        .Q(\bench_vout_reg[1] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [56]),
        .Q(\bench_vout_reg[1] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [57]),
        .Q(\bench_vout_reg[1] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [58]),
        .Q(\bench_vout_reg[1] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [59]),
        .Q(\bench_vout_reg[1] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [5]),
        .Q(\bench_vout_reg[1] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [60]),
        .Q(\bench_vout_reg[1] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [61]),
        .Q(\bench_vout_reg[1] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [62]),
        .Q(\bench_vout_reg[1] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [63]),
        .Q(\bench_vout_reg[1] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [64]),
        .Q(\bench_vout_reg[1] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [65]),
        .Q(\bench_vout_reg[1] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [66]),
        .Q(\bench_vout_reg[1] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [67]),
        .Q(\bench_vout_reg[1] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [68]),
        .Q(\bench_vout_reg[1] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [69]),
        .Q(\bench_vout_reg[1] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [6]),
        .Q(\bench_vout_reg[1] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [70]),
        .Q(\bench_vout_reg[1] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [71]),
        .Q(\bench_vout_reg[1] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [72]),
        .Q(\bench_vout_reg[1] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [73]),
        .Q(\bench_vout_reg[1] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [74]),
        .Q(\bench_vout_reg[1] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [75]),
        .Q(\bench_vout_reg[1] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [76]),
        .Q(\bench_vout_reg[1] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [77]),
        .Q(\bench_vout_reg[1] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [78]),
        .Q(\bench_vout_reg[1] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [79]),
        .Q(\bench_vout_reg[1] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [7]),
        .Q(\bench_vout_reg[1] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [80]),
        .Q(\bench_vout_reg[1] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [81]),
        .Q(\bench_vout_reg[1] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [82]),
        .Q(\bench_vout_reg[1] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [83]),
        .Q(\bench_vout_reg[1] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [84]),
        .Q(\bench_vout_reg[1] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [85]),
        .Q(\bench_vout_reg[1] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [86]),
        .Q(\bench_vout_reg[1] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [87]),
        .Q(\bench_vout_reg[1] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [88]),
        .Q(\bench_vout_reg[1] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [89]),
        .Q(\bench_vout_reg[1] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [8]),
        .Q(\bench_vout_reg[1] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [90]),
        .Q(\bench_vout_reg[1] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [91]),
        .Q(\bench_vout_reg[1] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [92]),
        .Q(\bench_vout_reg[1] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [93]),
        .Q(\bench_vout_reg[1] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [94]),
        .Q(\bench_vout_reg[1] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [95]),
        .Q(\bench_vout_reg[1] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [96]),
        .Q(\bench_vout_reg[1] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [97]),
        .Q(\bench_vout_reg[1] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [98]),
        .Q(\bench_vout_reg[1] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [99]),
        .Q(\bench_vout_reg[1] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[1].bench_vout_reg_reg[1][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[1] [9]),
        .Q(\bench_vout_reg[1] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng__2 \noise_circ_replica[1].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[1] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[1] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench__2 \noise_circ_replica[1].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[1] [24]),
        .g1006(\bench_vout[1] [7]),
        .g1008(\bench_v[1] [25]),
        .g1015(\bench_vout[1] [8]),
        .g1016(\bench_v[1] [26]),
        .g1017(\bench_vout[1] [9]),
        .g1080(\bench_v[1] [27]),
        .g1234(\bench_v[1] [28]),
        .g1246(\bench_vout[1] [10]),
        .g1553(\bench_v[1] [29]),
        .g1554(\bench_v[1] [30]),
        .g1724(\bench_vout[1] [11]),
        .g1783(\bench_vout[1] [12]),
        .g1798(\bench_vout[1] [13]),
        .g1804(\bench_vout[1] [14]),
        .g1810(\bench_vout[1] [15]),
        .g1817(\bench_vout[1] [16]),
        .g1824(\bench_vout[1] [17]),
        .g1829(\bench_vout[1] [18]),
        .g1870(\bench_vout[1] [19]),
        .g1871(\bench_vout[1] [20]),
        .g1894(\bench_vout[1] [21]),
        .g1911(\bench_vout[1] [22]),
        .g1944(\bench_vout[1] [23]),
        .g206(\bench_vout[1] [0]),
        .g2662(\bench_vout[1] [24]),
        .g2844(\bench_vout[1] [25]),
        .g2888(\bench_vout[1] [26]),
        .g291(\bench_vout[1] [1]),
        .g3077(\bench_vout[1] [27]),
        .g3096(\bench_vout[1] [28]),
        .g3130(\bench_vout[1] [29]),
        .g3159(\bench_vout[1] [30]),
        .g3191(\bench_vout[1] [31]),
        .g372(\bench_vout[1] [2]),
        .g3829(\bench_vout[1] [32]),
        .g3859(\bench_vout[1] [33]),
        .g3860(\bench_vout[1] [34]),
        .g4267(\bench_vout[1] [35]),
        .g43(\bench_v[1] [0]),
        .g4316(\bench_vout[1] [36]),
        .g4370(\bench_vout[1] [37]),
        .g4371(\bench_vout[1] [38]),
        .g4372(\bench_vout[1] [39]),
        .g4373(\bench_vout[1] [40]),
        .g453(\bench_vout[1] [3]),
        .g4655(\bench_vout[1] [41]),
        .g4657(\bench_vout[1] [42]),
        .g4660(\bench_vout[1] [43]),
        .g4661(\bench_vout[1] [44]),
        .g4663(\bench_vout[1] [45]),
        .g4664(\bench_vout[1] [46]),
        .g49(\bench_v[1] [1]),
        .g5143(\bench_vout[1] [47]),
        .g5164(\bench_vout[1] [48]),
        .g534(\bench_vout[1] [4]),
        .g5571(\bench_vout[1] [49]),
        .g5669(\bench_vout[1] [50]),
        .g5678(\bench_vout[1] [51]),
        .g5682(\bench_vout[1] [52]),
        .g5684(\bench_vout[1] [53]),
        .g5687(\bench_vout[1] [54]),
        .g5729(\bench_vout[1] [55]),
        .g594(\bench_vout[1] [5]),
        .g6207(\bench_vout[1] [56]),
        .g6212(\bench_vout[1] [57]),
        .g6223(\bench_vout[1] [58]),
        .g6236(\bench_vout[1] [59]),
        .g6269(\bench_vout[1] [60]),
        .g633(\bench_v[1] [2]),
        .g634(\bench_v[1] [3]),
        .g635(\bench_v[1] [4]),
        .g6425(\bench_vout[1] [61]),
        .g645(\bench_v[1] [5]),
        .g647(\bench_v[1] [6]),
        .g648(\bench_v[1] [7]),
        .g6648(\bench_vout[1] [62]),
        .g6653(\bench_vout[1] [63]),
        .g6675(\bench_vout[1] [64]),
        .g6849(\bench_vout[1] [65]),
        .g6850(\bench_vout[1] [66]),
        .g6895(\bench_vout[1] [67]),
        .g690(\bench_v[1] [8]),
        .g6909(\bench_vout[1] [68]),
        .g694(\bench_v[1] [9]),
        .g698(\bench_v[1] [10]),
        .g702(\bench_v[1] [11]),
        .g7048(\bench_vout[1] [69]),
        .g7063(\bench_vout[1] [70]),
        .g7103(\bench_vout[1] [71]),
        .g722(\bench_v[1] [12]),
        .g723(\bench_v[1] [13]),
        .g7283(\bench_vout[1] [72]),
        .g7284(\bench_vout[1] [73]),
        .g7285(\bench_vout[1] [74]),
        .g7286(\bench_vout[1] [75]),
        .g7287(\bench_vout[1] [76]),
        .g7288(\bench_vout[1] [77]),
        .g7289(\bench_vout[1] [78]),
        .g7290(\bench_vout[1] [79]),
        .g7291(\bench_vout[1] [80]),
        .g7292(\bench_vout[1] [81]),
        .g7293(\bench_vout[1] [82]),
        .g7294(\bench_vout[1] [83]),
        .g7295(\bench_vout[1] [84]),
        .g7298(\bench_vout[1] [85]),
        .g7423(\bench_vout[1] [86]),
        .g7424(\bench_vout[1] [87]),
        .g7425(\bench_vout[1] [88]),
        .g7474(\bench_vout[1] [89]),
        .g7504(\bench_vout[1] [90]),
        .g7505(\bench_vout[1] [91]),
        .g7506(\bench_vout[1] [92]),
        .g7507(\bench_vout[1] [93]),
        .g7508(\bench_vout[1] [94]),
        .g751(\bench_v[1] [14]),
        .g7514(\bench_vout[1] [95]),
        .g752(\bench_v[1] [15]),
        .g753(\bench_v[1] [16]),
        .g754(\bench_v[1] [17]),
        .g755(\bench_v[1] [18]),
        .g756(\bench_v[1] [19]),
        .g757(\bench_v[1] [20]),
        .g7729(\bench_vout[1] [96]),
        .g7730(\bench_vout[1] [97]),
        .g7731(\bench_vout[1] [98]),
        .g7732(\bench_vout[1] [99]),
        .g781(\bench_v[1] [21]),
        .g785(\bench_vout[1] [6]),
        .g8216(\bench_vout[1] [100]),
        .g8217(\bench_vout[1] [101]),
        .g8218(\bench_vout[1] [102]),
        .g8219(\bench_vout[1] [103]),
        .g8234(\bench_vout[1] [104]),
        .g8661(\bench_vout[1] [105]),
        .g8663(\bench_vout[1] [106]),
        .g8872(\bench_vout[1] [107]),
        .g8958(\bench_vout[1] [108]),
        .g9128(\bench_vout[1] [109]),
        .g9132(\bench_vout[1] [110]),
        .g9204(\bench_vout[1] [111]),
        .g9280(\bench_vout[1] [112]),
        .g9297(\bench_vout[1] [113]),
        .g9299(\bench_vout[1] [114]),
        .g9305(\bench_vout[1] [115]),
        .g9308(\bench_vout[1] [116]),
        .g9310(\bench_vout[1] [117]),
        .g9312(\bench_vout[1] [118]),
        .g9314(\bench_vout[1] [119]),
        .g9378(\bench_vout[1] [120]),
        .g941(\bench_v[1] [22]),
        .g962(\bench_v[1] [23]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [0]),
        .Q(\bench_vout_reg[2] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [100]),
        .Q(\bench_vout_reg[2] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [101]),
        .Q(\bench_vout_reg[2] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [102]),
        .Q(\bench_vout_reg[2] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [103]),
        .Q(\bench_vout_reg[2] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [104]),
        .Q(\bench_vout_reg[2] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [105]),
        .Q(\bench_vout_reg[2] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [106]),
        .Q(\bench_vout_reg[2] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [107]),
        .Q(\bench_vout_reg[2] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [108]),
        .Q(\bench_vout_reg[2] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [109]),
        .Q(\bench_vout_reg[2] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [10]),
        .Q(\bench_vout_reg[2] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [110]),
        .Q(\bench_vout_reg[2] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [111]),
        .Q(\bench_vout_reg[2] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [112]),
        .Q(\bench_vout_reg[2] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [113]),
        .Q(\bench_vout_reg[2] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [114]),
        .Q(\bench_vout_reg[2] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [115]),
        .Q(\bench_vout_reg[2] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [116]),
        .Q(\bench_vout_reg[2] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [117]),
        .Q(\bench_vout_reg[2] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [118]),
        .Q(\bench_vout_reg[2] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [119]),
        .Q(\bench_vout_reg[2] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [11]),
        .Q(\bench_vout_reg[2] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [120]),
        .Q(\bench_vout_reg[2] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [12]),
        .Q(\bench_vout_reg[2] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [13]),
        .Q(\bench_vout_reg[2] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [14]),
        .Q(\bench_vout_reg[2] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [15]),
        .Q(\bench_vout_reg[2] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [16]),
        .Q(\bench_vout_reg[2] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [17]),
        .Q(\bench_vout_reg[2] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [18]),
        .Q(\bench_vout_reg[2] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [19]),
        .Q(\bench_vout_reg[2] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [1]),
        .Q(\bench_vout_reg[2] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [20]),
        .Q(\bench_vout_reg[2] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [21]),
        .Q(\bench_vout_reg[2] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [22]),
        .Q(\bench_vout_reg[2] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [23]),
        .Q(\bench_vout_reg[2] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [24]),
        .Q(\bench_vout_reg[2] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [25]),
        .Q(\bench_vout_reg[2] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [26]),
        .Q(\bench_vout_reg[2] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [27]),
        .Q(\bench_vout_reg[2] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [28]),
        .Q(\bench_vout_reg[2] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [29]),
        .Q(\bench_vout_reg[2] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [2]),
        .Q(\bench_vout_reg[2] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [30]),
        .Q(\bench_vout_reg[2] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [31]),
        .Q(\bench_vout_reg[2] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [32]),
        .Q(\bench_vout_reg[2] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [33]),
        .Q(\bench_vout_reg[2] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [34]),
        .Q(\bench_vout_reg[2] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [35]),
        .Q(\bench_vout_reg[2] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [36]),
        .Q(\bench_vout_reg[2] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [37]),
        .Q(\bench_vout_reg[2] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [38]),
        .Q(\bench_vout_reg[2] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [39]),
        .Q(\bench_vout_reg[2] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [3]),
        .Q(\bench_vout_reg[2] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [40]),
        .Q(\bench_vout_reg[2] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [41]),
        .Q(\bench_vout_reg[2] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [42]),
        .Q(\bench_vout_reg[2] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [43]),
        .Q(\bench_vout_reg[2] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [44]),
        .Q(\bench_vout_reg[2] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [45]),
        .Q(\bench_vout_reg[2] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [46]),
        .Q(\bench_vout_reg[2] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [47]),
        .Q(\bench_vout_reg[2] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [48]),
        .Q(\bench_vout_reg[2] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [49]),
        .Q(\bench_vout_reg[2] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [4]),
        .Q(\bench_vout_reg[2] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [50]),
        .Q(\bench_vout_reg[2] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [51]),
        .Q(\bench_vout_reg[2] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [52]),
        .Q(\bench_vout_reg[2] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [53]),
        .Q(\bench_vout_reg[2] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [54]),
        .Q(\bench_vout_reg[2] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [55]),
        .Q(\bench_vout_reg[2] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [56]),
        .Q(\bench_vout_reg[2] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [57]),
        .Q(\bench_vout_reg[2] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [58]),
        .Q(\bench_vout_reg[2] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [59]),
        .Q(\bench_vout_reg[2] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [5]),
        .Q(\bench_vout_reg[2] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [60]),
        .Q(\bench_vout_reg[2] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [61]),
        .Q(\bench_vout_reg[2] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [62]),
        .Q(\bench_vout_reg[2] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [63]),
        .Q(\bench_vout_reg[2] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [64]),
        .Q(\bench_vout_reg[2] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [65]),
        .Q(\bench_vout_reg[2] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [66]),
        .Q(\bench_vout_reg[2] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [67]),
        .Q(\bench_vout_reg[2] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [68]),
        .Q(\bench_vout_reg[2] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [69]),
        .Q(\bench_vout_reg[2] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [6]),
        .Q(\bench_vout_reg[2] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [70]),
        .Q(\bench_vout_reg[2] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [71]),
        .Q(\bench_vout_reg[2] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [72]),
        .Q(\bench_vout_reg[2] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [73]),
        .Q(\bench_vout_reg[2] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [74]),
        .Q(\bench_vout_reg[2] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [75]),
        .Q(\bench_vout_reg[2] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [76]),
        .Q(\bench_vout_reg[2] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [77]),
        .Q(\bench_vout_reg[2] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [78]),
        .Q(\bench_vout_reg[2] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [79]),
        .Q(\bench_vout_reg[2] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [7]),
        .Q(\bench_vout_reg[2] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [80]),
        .Q(\bench_vout_reg[2] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [81]),
        .Q(\bench_vout_reg[2] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [82]),
        .Q(\bench_vout_reg[2] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [83]),
        .Q(\bench_vout_reg[2] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [84]),
        .Q(\bench_vout_reg[2] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [85]),
        .Q(\bench_vout_reg[2] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [86]),
        .Q(\bench_vout_reg[2] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [87]),
        .Q(\bench_vout_reg[2] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [88]),
        .Q(\bench_vout_reg[2] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [89]),
        .Q(\bench_vout_reg[2] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [8]),
        .Q(\bench_vout_reg[2] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [90]),
        .Q(\bench_vout_reg[2] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [91]),
        .Q(\bench_vout_reg[2] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [92]),
        .Q(\bench_vout_reg[2] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [93]),
        .Q(\bench_vout_reg[2] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [94]),
        .Q(\bench_vout_reg[2] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [95]),
        .Q(\bench_vout_reg[2] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [96]),
        .Q(\bench_vout_reg[2] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [97]),
        .Q(\bench_vout_reg[2] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [98]),
        .Q(\bench_vout_reg[2] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [99]),
        .Q(\bench_vout_reg[2] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[2].bench_vout_reg_reg[2][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[2] [9]),
        .Q(\bench_vout_reg[2] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng__3 \noise_circ_replica[2].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[2] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[2] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench__3 \noise_circ_replica[2].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[2] [24]),
        .g1006(\bench_vout[2] [7]),
        .g1008(\bench_v[2] [25]),
        .g1015(\bench_vout[2] [8]),
        .g1016(\bench_v[2] [26]),
        .g1017(\bench_vout[2] [9]),
        .g1080(\bench_v[2] [27]),
        .g1234(\bench_v[2] [28]),
        .g1246(\bench_vout[2] [10]),
        .g1553(\bench_v[2] [29]),
        .g1554(\bench_v[2] [30]),
        .g1724(\bench_vout[2] [11]),
        .g1783(\bench_vout[2] [12]),
        .g1798(\bench_vout[2] [13]),
        .g1804(\bench_vout[2] [14]),
        .g1810(\bench_vout[2] [15]),
        .g1817(\bench_vout[2] [16]),
        .g1824(\bench_vout[2] [17]),
        .g1829(\bench_vout[2] [18]),
        .g1870(\bench_vout[2] [19]),
        .g1871(\bench_vout[2] [20]),
        .g1894(\bench_vout[2] [21]),
        .g1911(\bench_vout[2] [22]),
        .g1944(\bench_vout[2] [23]),
        .g206(\bench_vout[2] [0]),
        .g2662(\bench_vout[2] [24]),
        .g2844(\bench_vout[2] [25]),
        .g2888(\bench_vout[2] [26]),
        .g291(\bench_vout[2] [1]),
        .g3077(\bench_vout[2] [27]),
        .g3096(\bench_vout[2] [28]),
        .g3130(\bench_vout[2] [29]),
        .g3159(\bench_vout[2] [30]),
        .g3191(\bench_vout[2] [31]),
        .g372(\bench_vout[2] [2]),
        .g3829(\bench_vout[2] [32]),
        .g3859(\bench_vout[2] [33]),
        .g3860(\bench_vout[2] [34]),
        .g4267(\bench_vout[2] [35]),
        .g43(\bench_v[2] [0]),
        .g4316(\bench_vout[2] [36]),
        .g4370(\bench_vout[2] [37]),
        .g4371(\bench_vout[2] [38]),
        .g4372(\bench_vout[2] [39]),
        .g4373(\bench_vout[2] [40]),
        .g453(\bench_vout[2] [3]),
        .g4655(\bench_vout[2] [41]),
        .g4657(\bench_vout[2] [42]),
        .g4660(\bench_vout[2] [43]),
        .g4661(\bench_vout[2] [44]),
        .g4663(\bench_vout[2] [45]),
        .g4664(\bench_vout[2] [46]),
        .g49(\bench_v[2] [1]),
        .g5143(\bench_vout[2] [47]),
        .g5164(\bench_vout[2] [48]),
        .g534(\bench_vout[2] [4]),
        .g5571(\bench_vout[2] [49]),
        .g5669(\bench_vout[2] [50]),
        .g5678(\bench_vout[2] [51]),
        .g5682(\bench_vout[2] [52]),
        .g5684(\bench_vout[2] [53]),
        .g5687(\bench_vout[2] [54]),
        .g5729(\bench_vout[2] [55]),
        .g594(\bench_vout[2] [5]),
        .g6207(\bench_vout[2] [56]),
        .g6212(\bench_vout[2] [57]),
        .g6223(\bench_vout[2] [58]),
        .g6236(\bench_vout[2] [59]),
        .g6269(\bench_vout[2] [60]),
        .g633(\bench_v[2] [2]),
        .g634(\bench_v[2] [3]),
        .g635(\bench_v[2] [4]),
        .g6425(\bench_vout[2] [61]),
        .g645(\bench_v[2] [5]),
        .g647(\bench_v[2] [6]),
        .g648(\bench_v[2] [7]),
        .g6648(\bench_vout[2] [62]),
        .g6653(\bench_vout[2] [63]),
        .g6675(\bench_vout[2] [64]),
        .g6849(\bench_vout[2] [65]),
        .g6850(\bench_vout[2] [66]),
        .g6895(\bench_vout[2] [67]),
        .g690(\bench_v[2] [8]),
        .g6909(\bench_vout[2] [68]),
        .g694(\bench_v[2] [9]),
        .g698(\bench_v[2] [10]),
        .g702(\bench_v[2] [11]),
        .g7048(\bench_vout[2] [69]),
        .g7063(\bench_vout[2] [70]),
        .g7103(\bench_vout[2] [71]),
        .g722(\bench_v[2] [12]),
        .g723(\bench_v[2] [13]),
        .g7283(\bench_vout[2] [72]),
        .g7284(\bench_vout[2] [73]),
        .g7285(\bench_vout[2] [74]),
        .g7286(\bench_vout[2] [75]),
        .g7287(\bench_vout[2] [76]),
        .g7288(\bench_vout[2] [77]),
        .g7289(\bench_vout[2] [78]),
        .g7290(\bench_vout[2] [79]),
        .g7291(\bench_vout[2] [80]),
        .g7292(\bench_vout[2] [81]),
        .g7293(\bench_vout[2] [82]),
        .g7294(\bench_vout[2] [83]),
        .g7295(\bench_vout[2] [84]),
        .g7298(\bench_vout[2] [85]),
        .g7423(\bench_vout[2] [86]),
        .g7424(\bench_vout[2] [87]),
        .g7425(\bench_vout[2] [88]),
        .g7474(\bench_vout[2] [89]),
        .g7504(\bench_vout[2] [90]),
        .g7505(\bench_vout[2] [91]),
        .g7506(\bench_vout[2] [92]),
        .g7507(\bench_vout[2] [93]),
        .g7508(\bench_vout[2] [94]),
        .g751(\bench_v[2] [14]),
        .g7514(\bench_vout[2] [95]),
        .g752(\bench_v[2] [15]),
        .g753(\bench_v[2] [16]),
        .g754(\bench_v[2] [17]),
        .g755(\bench_v[2] [18]),
        .g756(\bench_v[2] [19]),
        .g757(\bench_v[2] [20]),
        .g7729(\bench_vout[2] [96]),
        .g7730(\bench_vout[2] [97]),
        .g7731(\bench_vout[2] [98]),
        .g7732(\bench_vout[2] [99]),
        .g781(\bench_v[2] [21]),
        .g785(\bench_vout[2] [6]),
        .g8216(\bench_vout[2] [100]),
        .g8217(\bench_vout[2] [101]),
        .g8218(\bench_vout[2] [102]),
        .g8219(\bench_vout[2] [103]),
        .g8234(\bench_vout[2] [104]),
        .g8661(\bench_vout[2] [105]),
        .g8663(\bench_vout[2] [106]),
        .g8872(\bench_vout[2] [107]),
        .g8958(\bench_vout[2] [108]),
        .g9128(\bench_vout[2] [109]),
        .g9132(\bench_vout[2] [110]),
        .g9204(\bench_vout[2] [111]),
        .g9280(\bench_vout[2] [112]),
        .g9297(\bench_vout[2] [113]),
        .g9299(\bench_vout[2] [114]),
        .g9305(\bench_vout[2] [115]),
        .g9308(\bench_vout[2] [116]),
        .g9310(\bench_vout[2] [117]),
        .g9312(\bench_vout[2] [118]),
        .g9314(\bench_vout[2] [119]),
        .g9378(\bench_vout[2] [120]),
        .g941(\bench_v[2] [22]),
        .g962(\bench_v[2] [23]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [0]),
        .Q(\bench_vout_reg[3] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [100]),
        .Q(\bench_vout_reg[3] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [101]),
        .Q(\bench_vout_reg[3] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [102]),
        .Q(\bench_vout_reg[3] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [103]),
        .Q(\bench_vout_reg[3] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [104]),
        .Q(\bench_vout_reg[3] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [105]),
        .Q(\bench_vout_reg[3] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [106]),
        .Q(\bench_vout_reg[3] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [107]),
        .Q(\bench_vout_reg[3] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [108]),
        .Q(\bench_vout_reg[3] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [109]),
        .Q(\bench_vout_reg[3] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [10]),
        .Q(\bench_vout_reg[3] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [110]),
        .Q(\bench_vout_reg[3] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [111]),
        .Q(\bench_vout_reg[3] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [112]),
        .Q(\bench_vout_reg[3] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [113]),
        .Q(\bench_vout_reg[3] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [114]),
        .Q(\bench_vout_reg[3] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [115]),
        .Q(\bench_vout_reg[3] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [116]),
        .Q(\bench_vout_reg[3] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [117]),
        .Q(\bench_vout_reg[3] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [118]),
        .Q(\bench_vout_reg[3] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [119]),
        .Q(\bench_vout_reg[3] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [11]),
        .Q(\bench_vout_reg[3] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [120]),
        .Q(\bench_vout_reg[3] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [12]),
        .Q(\bench_vout_reg[3] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [13]),
        .Q(\bench_vout_reg[3] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [14]),
        .Q(\bench_vout_reg[3] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [15]),
        .Q(\bench_vout_reg[3] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [16]),
        .Q(\bench_vout_reg[3] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [17]),
        .Q(\bench_vout_reg[3] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [18]),
        .Q(\bench_vout_reg[3] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [19]),
        .Q(\bench_vout_reg[3] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [1]),
        .Q(\bench_vout_reg[3] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [20]),
        .Q(\bench_vout_reg[3] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [21]),
        .Q(\bench_vout_reg[3] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [22]),
        .Q(\bench_vout_reg[3] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [23]),
        .Q(\bench_vout_reg[3] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [24]),
        .Q(\bench_vout_reg[3] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [25]),
        .Q(\bench_vout_reg[3] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [26]),
        .Q(\bench_vout_reg[3] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [27]),
        .Q(\bench_vout_reg[3] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [28]),
        .Q(\bench_vout_reg[3] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [29]),
        .Q(\bench_vout_reg[3] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [2]),
        .Q(\bench_vout_reg[3] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [30]),
        .Q(\bench_vout_reg[3] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [31]),
        .Q(\bench_vout_reg[3] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [32]),
        .Q(\bench_vout_reg[3] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [33]),
        .Q(\bench_vout_reg[3] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [34]),
        .Q(\bench_vout_reg[3] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [35]),
        .Q(\bench_vout_reg[3] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [36]),
        .Q(\bench_vout_reg[3] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [37]),
        .Q(\bench_vout_reg[3] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [38]),
        .Q(\bench_vout_reg[3] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [39]),
        .Q(\bench_vout_reg[3] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [3]),
        .Q(\bench_vout_reg[3] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [40]),
        .Q(\bench_vout_reg[3] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [41]),
        .Q(\bench_vout_reg[3] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [42]),
        .Q(\bench_vout_reg[3] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [43]),
        .Q(\bench_vout_reg[3] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [44]),
        .Q(\bench_vout_reg[3] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [45]),
        .Q(\bench_vout_reg[3] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [46]),
        .Q(\bench_vout_reg[3] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [47]),
        .Q(\bench_vout_reg[3] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [48]),
        .Q(\bench_vout_reg[3] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [49]),
        .Q(\bench_vout_reg[3] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [4]),
        .Q(\bench_vout_reg[3] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [50]),
        .Q(\bench_vout_reg[3] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [51]),
        .Q(\bench_vout_reg[3] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [52]),
        .Q(\bench_vout_reg[3] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [53]),
        .Q(\bench_vout_reg[3] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [54]),
        .Q(\bench_vout_reg[3] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [55]),
        .Q(\bench_vout_reg[3] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [56]),
        .Q(\bench_vout_reg[3] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [57]),
        .Q(\bench_vout_reg[3] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [58]),
        .Q(\bench_vout_reg[3] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [59]),
        .Q(\bench_vout_reg[3] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [5]),
        .Q(\bench_vout_reg[3] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [60]),
        .Q(\bench_vout_reg[3] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [61]),
        .Q(\bench_vout_reg[3] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [62]),
        .Q(\bench_vout_reg[3] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [63]),
        .Q(\bench_vout_reg[3] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [64]),
        .Q(\bench_vout_reg[3] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [65]),
        .Q(\bench_vout_reg[3] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [66]),
        .Q(\bench_vout_reg[3] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [67]),
        .Q(\bench_vout_reg[3] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [68]),
        .Q(\bench_vout_reg[3] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [69]),
        .Q(\bench_vout_reg[3] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [6]),
        .Q(\bench_vout_reg[3] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [70]),
        .Q(\bench_vout_reg[3] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [71]),
        .Q(\bench_vout_reg[3] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [72]),
        .Q(\bench_vout_reg[3] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [73]),
        .Q(\bench_vout_reg[3] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [74]),
        .Q(\bench_vout_reg[3] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [75]),
        .Q(\bench_vout_reg[3] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [76]),
        .Q(\bench_vout_reg[3] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [77]),
        .Q(\bench_vout_reg[3] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [78]),
        .Q(\bench_vout_reg[3] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [79]),
        .Q(\bench_vout_reg[3] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [7]),
        .Q(\bench_vout_reg[3] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [80]),
        .Q(\bench_vout_reg[3] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [81]),
        .Q(\bench_vout_reg[3] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [82]),
        .Q(\bench_vout_reg[3] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [83]),
        .Q(\bench_vout_reg[3] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [84]),
        .Q(\bench_vout_reg[3] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [85]),
        .Q(\bench_vout_reg[3] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [86]),
        .Q(\bench_vout_reg[3] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [87]),
        .Q(\bench_vout_reg[3] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [88]),
        .Q(\bench_vout_reg[3] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [89]),
        .Q(\bench_vout_reg[3] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [8]),
        .Q(\bench_vout_reg[3] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [90]),
        .Q(\bench_vout_reg[3] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [91]),
        .Q(\bench_vout_reg[3] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [92]),
        .Q(\bench_vout_reg[3] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [93]),
        .Q(\bench_vout_reg[3] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [94]),
        .Q(\bench_vout_reg[3] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [95]),
        .Q(\bench_vout_reg[3] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [96]),
        .Q(\bench_vout_reg[3] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [97]),
        .Q(\bench_vout_reg[3] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [98]),
        .Q(\bench_vout_reg[3] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [99]),
        .Q(\bench_vout_reg[3] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[3].bench_vout_reg_reg[3][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[3] [9]),
        .Q(\bench_vout_reg[3] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng__4 \noise_circ_replica[3].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[3] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[3] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench__4 \noise_circ_replica[3].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[3] [24]),
        .g1006(\bench_vout[3] [7]),
        .g1008(\bench_v[3] [25]),
        .g1015(\bench_vout[3] [8]),
        .g1016(\bench_v[3] [26]),
        .g1017(\bench_vout[3] [9]),
        .g1080(\bench_v[3] [27]),
        .g1234(\bench_v[3] [28]),
        .g1246(\bench_vout[3] [10]),
        .g1553(\bench_v[3] [29]),
        .g1554(\bench_v[3] [30]),
        .g1724(\bench_vout[3] [11]),
        .g1783(\bench_vout[3] [12]),
        .g1798(\bench_vout[3] [13]),
        .g1804(\bench_vout[3] [14]),
        .g1810(\bench_vout[3] [15]),
        .g1817(\bench_vout[3] [16]),
        .g1824(\bench_vout[3] [17]),
        .g1829(\bench_vout[3] [18]),
        .g1870(\bench_vout[3] [19]),
        .g1871(\bench_vout[3] [20]),
        .g1894(\bench_vout[3] [21]),
        .g1911(\bench_vout[3] [22]),
        .g1944(\bench_vout[3] [23]),
        .g206(\bench_vout[3] [0]),
        .g2662(\bench_vout[3] [24]),
        .g2844(\bench_vout[3] [25]),
        .g2888(\bench_vout[3] [26]),
        .g291(\bench_vout[3] [1]),
        .g3077(\bench_vout[3] [27]),
        .g3096(\bench_vout[3] [28]),
        .g3130(\bench_vout[3] [29]),
        .g3159(\bench_vout[3] [30]),
        .g3191(\bench_vout[3] [31]),
        .g372(\bench_vout[3] [2]),
        .g3829(\bench_vout[3] [32]),
        .g3859(\bench_vout[3] [33]),
        .g3860(\bench_vout[3] [34]),
        .g4267(\bench_vout[3] [35]),
        .g43(\bench_v[3] [0]),
        .g4316(\bench_vout[3] [36]),
        .g4370(\bench_vout[3] [37]),
        .g4371(\bench_vout[3] [38]),
        .g4372(\bench_vout[3] [39]),
        .g4373(\bench_vout[3] [40]),
        .g453(\bench_vout[3] [3]),
        .g4655(\bench_vout[3] [41]),
        .g4657(\bench_vout[3] [42]),
        .g4660(\bench_vout[3] [43]),
        .g4661(\bench_vout[3] [44]),
        .g4663(\bench_vout[3] [45]),
        .g4664(\bench_vout[3] [46]),
        .g49(\bench_v[3] [1]),
        .g5143(\bench_vout[3] [47]),
        .g5164(\bench_vout[3] [48]),
        .g534(\bench_vout[3] [4]),
        .g5571(\bench_vout[3] [49]),
        .g5669(\bench_vout[3] [50]),
        .g5678(\bench_vout[3] [51]),
        .g5682(\bench_vout[3] [52]),
        .g5684(\bench_vout[3] [53]),
        .g5687(\bench_vout[3] [54]),
        .g5729(\bench_vout[3] [55]),
        .g594(\bench_vout[3] [5]),
        .g6207(\bench_vout[3] [56]),
        .g6212(\bench_vout[3] [57]),
        .g6223(\bench_vout[3] [58]),
        .g6236(\bench_vout[3] [59]),
        .g6269(\bench_vout[3] [60]),
        .g633(\bench_v[3] [2]),
        .g634(\bench_v[3] [3]),
        .g635(\bench_v[3] [4]),
        .g6425(\bench_vout[3] [61]),
        .g645(\bench_v[3] [5]),
        .g647(\bench_v[3] [6]),
        .g648(\bench_v[3] [7]),
        .g6648(\bench_vout[3] [62]),
        .g6653(\bench_vout[3] [63]),
        .g6675(\bench_vout[3] [64]),
        .g6849(\bench_vout[3] [65]),
        .g6850(\bench_vout[3] [66]),
        .g6895(\bench_vout[3] [67]),
        .g690(\bench_v[3] [8]),
        .g6909(\bench_vout[3] [68]),
        .g694(\bench_v[3] [9]),
        .g698(\bench_v[3] [10]),
        .g702(\bench_v[3] [11]),
        .g7048(\bench_vout[3] [69]),
        .g7063(\bench_vout[3] [70]),
        .g7103(\bench_vout[3] [71]),
        .g722(\bench_v[3] [12]),
        .g723(\bench_v[3] [13]),
        .g7283(\bench_vout[3] [72]),
        .g7284(\bench_vout[3] [73]),
        .g7285(\bench_vout[3] [74]),
        .g7286(\bench_vout[3] [75]),
        .g7287(\bench_vout[3] [76]),
        .g7288(\bench_vout[3] [77]),
        .g7289(\bench_vout[3] [78]),
        .g7290(\bench_vout[3] [79]),
        .g7291(\bench_vout[3] [80]),
        .g7292(\bench_vout[3] [81]),
        .g7293(\bench_vout[3] [82]),
        .g7294(\bench_vout[3] [83]),
        .g7295(\bench_vout[3] [84]),
        .g7298(\bench_vout[3] [85]),
        .g7423(\bench_vout[3] [86]),
        .g7424(\bench_vout[3] [87]),
        .g7425(\bench_vout[3] [88]),
        .g7474(\bench_vout[3] [89]),
        .g7504(\bench_vout[3] [90]),
        .g7505(\bench_vout[3] [91]),
        .g7506(\bench_vout[3] [92]),
        .g7507(\bench_vout[3] [93]),
        .g7508(\bench_vout[3] [94]),
        .g751(\bench_v[3] [14]),
        .g7514(\bench_vout[3] [95]),
        .g752(\bench_v[3] [15]),
        .g753(\bench_v[3] [16]),
        .g754(\bench_v[3] [17]),
        .g755(\bench_v[3] [18]),
        .g756(\bench_v[3] [19]),
        .g757(\bench_v[3] [20]),
        .g7729(\bench_vout[3] [96]),
        .g7730(\bench_vout[3] [97]),
        .g7731(\bench_vout[3] [98]),
        .g7732(\bench_vout[3] [99]),
        .g781(\bench_v[3] [21]),
        .g785(\bench_vout[3] [6]),
        .g8216(\bench_vout[3] [100]),
        .g8217(\bench_vout[3] [101]),
        .g8218(\bench_vout[3] [102]),
        .g8219(\bench_vout[3] [103]),
        .g8234(\bench_vout[3] [104]),
        .g8661(\bench_vout[3] [105]),
        .g8663(\bench_vout[3] [106]),
        .g8872(\bench_vout[3] [107]),
        .g8958(\bench_vout[3] [108]),
        .g9128(\bench_vout[3] [109]),
        .g9132(\bench_vout[3] [110]),
        .g9204(\bench_vout[3] [111]),
        .g9280(\bench_vout[3] [112]),
        .g9297(\bench_vout[3] [113]),
        .g9299(\bench_vout[3] [114]),
        .g9305(\bench_vout[3] [115]),
        .g9308(\bench_vout[3] [116]),
        .g9310(\bench_vout[3] [117]),
        .g9312(\bench_vout[3] [118]),
        .g9314(\bench_vout[3] [119]),
        .g9378(\bench_vout[3] [120]),
        .g941(\bench_v[3] [22]),
        .g962(\bench_v[3] [23]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [0]),
        .Q(\bench_vout_reg[4] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [100]),
        .Q(\bench_vout_reg[4] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [101]),
        .Q(\bench_vout_reg[4] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [102]),
        .Q(\bench_vout_reg[4] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [103]),
        .Q(\bench_vout_reg[4] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [104]),
        .Q(\bench_vout_reg[4] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [105]),
        .Q(\bench_vout_reg[4] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [106]),
        .Q(\bench_vout_reg[4] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [107]),
        .Q(\bench_vout_reg[4] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [108]),
        .Q(\bench_vout_reg[4] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [109]),
        .Q(\bench_vout_reg[4] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [10]),
        .Q(\bench_vout_reg[4] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [110]),
        .Q(\bench_vout_reg[4] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [111]),
        .Q(\bench_vout_reg[4] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [112]),
        .Q(\bench_vout_reg[4] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [113]),
        .Q(\bench_vout_reg[4] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [114]),
        .Q(\bench_vout_reg[4] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [115]),
        .Q(\bench_vout_reg[4] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [116]),
        .Q(\bench_vout_reg[4] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [117]),
        .Q(\bench_vout_reg[4] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [118]),
        .Q(\bench_vout_reg[4] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [119]),
        .Q(\bench_vout_reg[4] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [11]),
        .Q(\bench_vout_reg[4] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [120]),
        .Q(\bench_vout_reg[4] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [12]),
        .Q(\bench_vout_reg[4] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [13]),
        .Q(\bench_vout_reg[4] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [14]),
        .Q(\bench_vout_reg[4] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [15]),
        .Q(\bench_vout_reg[4] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [16]),
        .Q(\bench_vout_reg[4] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [17]),
        .Q(\bench_vout_reg[4] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [18]),
        .Q(\bench_vout_reg[4] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [19]),
        .Q(\bench_vout_reg[4] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [1]),
        .Q(\bench_vout_reg[4] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [20]),
        .Q(\bench_vout_reg[4] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [21]),
        .Q(\bench_vout_reg[4] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [22]),
        .Q(\bench_vout_reg[4] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [23]),
        .Q(\bench_vout_reg[4] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [24]),
        .Q(\bench_vout_reg[4] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [25]),
        .Q(\bench_vout_reg[4] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [26]),
        .Q(\bench_vout_reg[4] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [27]),
        .Q(\bench_vout_reg[4] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [28]),
        .Q(\bench_vout_reg[4] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [29]),
        .Q(\bench_vout_reg[4] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [2]),
        .Q(\bench_vout_reg[4] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [30]),
        .Q(\bench_vout_reg[4] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [31]),
        .Q(\bench_vout_reg[4] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [32]),
        .Q(\bench_vout_reg[4] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [33]),
        .Q(\bench_vout_reg[4] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [34]),
        .Q(\bench_vout_reg[4] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [35]),
        .Q(\bench_vout_reg[4] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [36]),
        .Q(\bench_vout_reg[4] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [37]),
        .Q(\bench_vout_reg[4] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [38]),
        .Q(\bench_vout_reg[4] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [39]),
        .Q(\bench_vout_reg[4] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [3]),
        .Q(\bench_vout_reg[4] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [40]),
        .Q(\bench_vout_reg[4] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [41]),
        .Q(\bench_vout_reg[4] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [42]),
        .Q(\bench_vout_reg[4] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [43]),
        .Q(\bench_vout_reg[4] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [44]),
        .Q(\bench_vout_reg[4] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [45]),
        .Q(\bench_vout_reg[4] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [46]),
        .Q(\bench_vout_reg[4] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [47]),
        .Q(\bench_vout_reg[4] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [48]),
        .Q(\bench_vout_reg[4] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [49]),
        .Q(\bench_vout_reg[4] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [4]),
        .Q(\bench_vout_reg[4] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [50]),
        .Q(\bench_vout_reg[4] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [51]),
        .Q(\bench_vout_reg[4] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [52]),
        .Q(\bench_vout_reg[4] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [53]),
        .Q(\bench_vout_reg[4] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [54]),
        .Q(\bench_vout_reg[4] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [55]),
        .Q(\bench_vout_reg[4] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [56]),
        .Q(\bench_vout_reg[4] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [57]),
        .Q(\bench_vout_reg[4] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [58]),
        .Q(\bench_vout_reg[4] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [59]),
        .Q(\bench_vout_reg[4] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [5]),
        .Q(\bench_vout_reg[4] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [60]),
        .Q(\bench_vout_reg[4] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [61]),
        .Q(\bench_vout_reg[4] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [62]),
        .Q(\bench_vout_reg[4] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [63]),
        .Q(\bench_vout_reg[4] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [64]),
        .Q(\bench_vout_reg[4] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [65]),
        .Q(\bench_vout_reg[4] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [66]),
        .Q(\bench_vout_reg[4] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [67]),
        .Q(\bench_vout_reg[4] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [68]),
        .Q(\bench_vout_reg[4] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [69]),
        .Q(\bench_vout_reg[4] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [6]),
        .Q(\bench_vout_reg[4] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [70]),
        .Q(\bench_vout_reg[4] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [71]),
        .Q(\bench_vout_reg[4] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [72]),
        .Q(\bench_vout_reg[4] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [73]),
        .Q(\bench_vout_reg[4] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [74]),
        .Q(\bench_vout_reg[4] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [75]),
        .Q(\bench_vout_reg[4] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [76]),
        .Q(\bench_vout_reg[4] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [77]),
        .Q(\bench_vout_reg[4] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [78]),
        .Q(\bench_vout_reg[4] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [79]),
        .Q(\bench_vout_reg[4] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [7]),
        .Q(\bench_vout_reg[4] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [80]),
        .Q(\bench_vout_reg[4] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [81]),
        .Q(\bench_vout_reg[4] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [82]),
        .Q(\bench_vout_reg[4] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [83]),
        .Q(\bench_vout_reg[4] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [84]),
        .Q(\bench_vout_reg[4] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [85]),
        .Q(\bench_vout_reg[4] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [86]),
        .Q(\bench_vout_reg[4] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [87]),
        .Q(\bench_vout_reg[4] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [88]),
        .Q(\bench_vout_reg[4] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [89]),
        .Q(\bench_vout_reg[4] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [8]),
        .Q(\bench_vout_reg[4] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [90]),
        .Q(\bench_vout_reg[4] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [91]),
        .Q(\bench_vout_reg[4] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [92]),
        .Q(\bench_vout_reg[4] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [93]),
        .Q(\bench_vout_reg[4] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [94]),
        .Q(\bench_vout_reg[4] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [95]),
        .Q(\bench_vout_reg[4] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [96]),
        .Q(\bench_vout_reg[4] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [97]),
        .Q(\bench_vout_reg[4] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [98]),
        .Q(\bench_vout_reg[4] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [99]),
        .Q(\bench_vout_reg[4] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[4].bench_vout_reg_reg[4][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[4] [9]),
        .Q(\bench_vout_reg[4] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng__5 \noise_circ_replica[4].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[4] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[4] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench__5 \noise_circ_replica[4].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[4] [24]),
        .g1006(\bench_vout[4] [7]),
        .g1008(\bench_v[4] [25]),
        .g1015(\bench_vout[4] [8]),
        .g1016(\bench_v[4] [26]),
        .g1017(\bench_vout[4] [9]),
        .g1080(\bench_v[4] [27]),
        .g1234(\bench_v[4] [28]),
        .g1246(\bench_vout[4] [10]),
        .g1553(\bench_v[4] [29]),
        .g1554(\bench_v[4] [30]),
        .g1724(\bench_vout[4] [11]),
        .g1783(\bench_vout[4] [12]),
        .g1798(\bench_vout[4] [13]),
        .g1804(\bench_vout[4] [14]),
        .g1810(\bench_vout[4] [15]),
        .g1817(\bench_vout[4] [16]),
        .g1824(\bench_vout[4] [17]),
        .g1829(\bench_vout[4] [18]),
        .g1870(\bench_vout[4] [19]),
        .g1871(\bench_vout[4] [20]),
        .g1894(\bench_vout[4] [21]),
        .g1911(\bench_vout[4] [22]),
        .g1944(\bench_vout[4] [23]),
        .g206(\bench_vout[4] [0]),
        .g2662(\bench_vout[4] [24]),
        .g2844(\bench_vout[4] [25]),
        .g2888(\bench_vout[4] [26]),
        .g291(\bench_vout[4] [1]),
        .g3077(\bench_vout[4] [27]),
        .g3096(\bench_vout[4] [28]),
        .g3130(\bench_vout[4] [29]),
        .g3159(\bench_vout[4] [30]),
        .g3191(\bench_vout[4] [31]),
        .g372(\bench_vout[4] [2]),
        .g3829(\bench_vout[4] [32]),
        .g3859(\bench_vout[4] [33]),
        .g3860(\bench_vout[4] [34]),
        .g4267(\bench_vout[4] [35]),
        .g43(\bench_v[4] [0]),
        .g4316(\bench_vout[4] [36]),
        .g4370(\bench_vout[4] [37]),
        .g4371(\bench_vout[4] [38]),
        .g4372(\bench_vout[4] [39]),
        .g4373(\bench_vout[4] [40]),
        .g453(\bench_vout[4] [3]),
        .g4655(\bench_vout[4] [41]),
        .g4657(\bench_vout[4] [42]),
        .g4660(\bench_vout[4] [43]),
        .g4661(\bench_vout[4] [44]),
        .g4663(\bench_vout[4] [45]),
        .g4664(\bench_vout[4] [46]),
        .g49(\bench_v[4] [1]),
        .g5143(\bench_vout[4] [47]),
        .g5164(\bench_vout[4] [48]),
        .g534(\bench_vout[4] [4]),
        .g5571(\bench_vout[4] [49]),
        .g5669(\bench_vout[4] [50]),
        .g5678(\bench_vout[4] [51]),
        .g5682(\bench_vout[4] [52]),
        .g5684(\bench_vout[4] [53]),
        .g5687(\bench_vout[4] [54]),
        .g5729(\bench_vout[4] [55]),
        .g594(\bench_vout[4] [5]),
        .g6207(\bench_vout[4] [56]),
        .g6212(\bench_vout[4] [57]),
        .g6223(\bench_vout[4] [58]),
        .g6236(\bench_vout[4] [59]),
        .g6269(\bench_vout[4] [60]),
        .g633(\bench_v[4] [2]),
        .g634(\bench_v[4] [3]),
        .g635(\bench_v[4] [4]),
        .g6425(\bench_vout[4] [61]),
        .g645(\bench_v[4] [5]),
        .g647(\bench_v[4] [6]),
        .g648(\bench_v[4] [7]),
        .g6648(\bench_vout[4] [62]),
        .g6653(\bench_vout[4] [63]),
        .g6675(\bench_vout[4] [64]),
        .g6849(\bench_vout[4] [65]),
        .g6850(\bench_vout[4] [66]),
        .g6895(\bench_vout[4] [67]),
        .g690(\bench_v[4] [8]),
        .g6909(\bench_vout[4] [68]),
        .g694(\bench_v[4] [9]),
        .g698(\bench_v[4] [10]),
        .g702(\bench_v[4] [11]),
        .g7048(\bench_vout[4] [69]),
        .g7063(\bench_vout[4] [70]),
        .g7103(\bench_vout[4] [71]),
        .g722(\bench_v[4] [12]),
        .g723(\bench_v[4] [13]),
        .g7283(\bench_vout[4] [72]),
        .g7284(\bench_vout[4] [73]),
        .g7285(\bench_vout[4] [74]),
        .g7286(\bench_vout[4] [75]),
        .g7287(\bench_vout[4] [76]),
        .g7288(\bench_vout[4] [77]),
        .g7289(\bench_vout[4] [78]),
        .g7290(\bench_vout[4] [79]),
        .g7291(\bench_vout[4] [80]),
        .g7292(\bench_vout[4] [81]),
        .g7293(\bench_vout[4] [82]),
        .g7294(\bench_vout[4] [83]),
        .g7295(\bench_vout[4] [84]),
        .g7298(\bench_vout[4] [85]),
        .g7423(\bench_vout[4] [86]),
        .g7424(\bench_vout[4] [87]),
        .g7425(\bench_vout[4] [88]),
        .g7474(\bench_vout[4] [89]),
        .g7504(\bench_vout[4] [90]),
        .g7505(\bench_vout[4] [91]),
        .g7506(\bench_vout[4] [92]),
        .g7507(\bench_vout[4] [93]),
        .g7508(\bench_vout[4] [94]),
        .g751(\bench_v[4] [14]),
        .g7514(\bench_vout[4] [95]),
        .g752(\bench_v[4] [15]),
        .g753(\bench_v[4] [16]),
        .g754(\bench_v[4] [17]),
        .g755(\bench_v[4] [18]),
        .g756(\bench_v[4] [19]),
        .g757(\bench_v[4] [20]),
        .g7729(\bench_vout[4] [96]),
        .g7730(\bench_vout[4] [97]),
        .g7731(\bench_vout[4] [98]),
        .g7732(\bench_vout[4] [99]),
        .g781(\bench_v[4] [21]),
        .g785(\bench_vout[4] [6]),
        .g8216(\bench_vout[4] [100]),
        .g8217(\bench_vout[4] [101]),
        .g8218(\bench_vout[4] [102]),
        .g8219(\bench_vout[4] [103]),
        .g8234(\bench_vout[4] [104]),
        .g8661(\bench_vout[4] [105]),
        .g8663(\bench_vout[4] [106]),
        .g8872(\bench_vout[4] [107]),
        .g8958(\bench_vout[4] [108]),
        .g9128(\bench_vout[4] [109]),
        .g9132(\bench_vout[4] [110]),
        .g9204(\bench_vout[4] [111]),
        .g9280(\bench_vout[4] [112]),
        .g9297(\bench_vout[4] [113]),
        .g9299(\bench_vout[4] [114]),
        .g9305(\bench_vout[4] [115]),
        .g9308(\bench_vout[4] [116]),
        .g9310(\bench_vout[4] [117]),
        .g9312(\bench_vout[4] [118]),
        .g9314(\bench_vout[4] [119]),
        .g9378(\bench_vout[4] [120]),
        .g941(\bench_v[4] [22]),
        .g962(\bench_v[4] [23]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [0]),
        .Q(\bench_vout_reg[5] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [100]),
        .Q(\bench_vout_reg[5] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [101]),
        .Q(\bench_vout_reg[5] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [102]),
        .Q(\bench_vout_reg[5] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [103]),
        .Q(\bench_vout_reg[5] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [104]),
        .Q(\bench_vout_reg[5] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [105]),
        .Q(\bench_vout_reg[5] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [106]),
        .Q(\bench_vout_reg[5] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [107]),
        .Q(\bench_vout_reg[5] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [108]),
        .Q(\bench_vout_reg[5] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [109]),
        .Q(\bench_vout_reg[5] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [10]),
        .Q(\bench_vout_reg[5] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [110]),
        .Q(\bench_vout_reg[5] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [111]),
        .Q(\bench_vout_reg[5] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [112]),
        .Q(\bench_vout_reg[5] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [113]),
        .Q(\bench_vout_reg[5] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [114]),
        .Q(\bench_vout_reg[5] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [115]),
        .Q(\bench_vout_reg[5] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [116]),
        .Q(\bench_vout_reg[5] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [117]),
        .Q(\bench_vout_reg[5] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [118]),
        .Q(\bench_vout_reg[5] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [119]),
        .Q(\bench_vout_reg[5] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [11]),
        .Q(\bench_vout_reg[5] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [120]),
        .Q(\bench_vout_reg[5] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [12]),
        .Q(\bench_vout_reg[5] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [13]),
        .Q(\bench_vout_reg[5] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [14]),
        .Q(\bench_vout_reg[5] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [15]),
        .Q(\bench_vout_reg[5] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [16]),
        .Q(\bench_vout_reg[5] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [17]),
        .Q(\bench_vout_reg[5] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [18]),
        .Q(\bench_vout_reg[5] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [19]),
        .Q(\bench_vout_reg[5] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [1]),
        .Q(\bench_vout_reg[5] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [20]),
        .Q(\bench_vout_reg[5] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [21]),
        .Q(\bench_vout_reg[5] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [22]),
        .Q(\bench_vout_reg[5] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [23]),
        .Q(\bench_vout_reg[5] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [24]),
        .Q(\bench_vout_reg[5] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [25]),
        .Q(\bench_vout_reg[5] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [26]),
        .Q(\bench_vout_reg[5] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [27]),
        .Q(\bench_vout_reg[5] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [28]),
        .Q(\bench_vout_reg[5] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [29]),
        .Q(\bench_vout_reg[5] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [2]),
        .Q(\bench_vout_reg[5] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [30]),
        .Q(\bench_vout_reg[5] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [31]),
        .Q(\bench_vout_reg[5] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [32]),
        .Q(\bench_vout_reg[5] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [33]),
        .Q(\bench_vout_reg[5] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [34]),
        .Q(\bench_vout_reg[5] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [35]),
        .Q(\bench_vout_reg[5] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [36]),
        .Q(\bench_vout_reg[5] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [37]),
        .Q(\bench_vout_reg[5] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [38]),
        .Q(\bench_vout_reg[5] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [39]),
        .Q(\bench_vout_reg[5] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [3]),
        .Q(\bench_vout_reg[5] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [40]),
        .Q(\bench_vout_reg[5] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [41]),
        .Q(\bench_vout_reg[5] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [42]),
        .Q(\bench_vout_reg[5] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [43]),
        .Q(\bench_vout_reg[5] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [44]),
        .Q(\bench_vout_reg[5] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [45]),
        .Q(\bench_vout_reg[5] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [46]),
        .Q(\bench_vout_reg[5] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [47]),
        .Q(\bench_vout_reg[5] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [48]),
        .Q(\bench_vout_reg[5] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [49]),
        .Q(\bench_vout_reg[5] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [4]),
        .Q(\bench_vout_reg[5] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [50]),
        .Q(\bench_vout_reg[5] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [51]),
        .Q(\bench_vout_reg[5] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [52]),
        .Q(\bench_vout_reg[5] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [53]),
        .Q(\bench_vout_reg[5] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [54]),
        .Q(\bench_vout_reg[5] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [55]),
        .Q(\bench_vout_reg[5] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [56]),
        .Q(\bench_vout_reg[5] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [57]),
        .Q(\bench_vout_reg[5] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [58]),
        .Q(\bench_vout_reg[5] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [59]),
        .Q(\bench_vout_reg[5] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [5]),
        .Q(\bench_vout_reg[5] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [60]),
        .Q(\bench_vout_reg[5] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [61]),
        .Q(\bench_vout_reg[5] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [62]),
        .Q(\bench_vout_reg[5] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [63]),
        .Q(\bench_vout_reg[5] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [64]),
        .Q(\bench_vout_reg[5] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [65]),
        .Q(\bench_vout_reg[5] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [66]),
        .Q(\bench_vout_reg[5] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [67]),
        .Q(\bench_vout_reg[5] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [68]),
        .Q(\bench_vout_reg[5] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [69]),
        .Q(\bench_vout_reg[5] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [6]),
        .Q(\bench_vout_reg[5] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [70]),
        .Q(\bench_vout_reg[5] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [71]),
        .Q(\bench_vout_reg[5] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [72]),
        .Q(\bench_vout_reg[5] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [73]),
        .Q(\bench_vout_reg[5] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [74]),
        .Q(\bench_vout_reg[5] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [75]),
        .Q(\bench_vout_reg[5] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [76]),
        .Q(\bench_vout_reg[5] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [77]),
        .Q(\bench_vout_reg[5] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [78]),
        .Q(\bench_vout_reg[5] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [79]),
        .Q(\bench_vout_reg[5] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [7]),
        .Q(\bench_vout_reg[5] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [80]),
        .Q(\bench_vout_reg[5] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [81]),
        .Q(\bench_vout_reg[5] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [82]),
        .Q(\bench_vout_reg[5] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [83]),
        .Q(\bench_vout_reg[5] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [84]),
        .Q(\bench_vout_reg[5] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [85]),
        .Q(\bench_vout_reg[5] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [86]),
        .Q(\bench_vout_reg[5] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [87]),
        .Q(\bench_vout_reg[5] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [88]),
        .Q(\bench_vout_reg[5] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [89]),
        .Q(\bench_vout_reg[5] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [8]),
        .Q(\bench_vout_reg[5] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [90]),
        .Q(\bench_vout_reg[5] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [91]),
        .Q(\bench_vout_reg[5] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [92]),
        .Q(\bench_vout_reg[5] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [93]),
        .Q(\bench_vout_reg[5] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [94]),
        .Q(\bench_vout_reg[5] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [95]),
        .Q(\bench_vout_reg[5] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [96]),
        .Q(\bench_vout_reg[5] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [97]),
        .Q(\bench_vout_reg[5] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [98]),
        .Q(\bench_vout_reg[5] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [99]),
        .Q(\bench_vout_reg[5] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[5].bench_vout_reg_reg[5][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[5] [9]),
        .Q(\bench_vout_reg[5] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng__6 \noise_circ_replica[5].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[5] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[5] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench__6 \noise_circ_replica[5].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[5] [24]),
        .g1006(\bench_vout[5] [7]),
        .g1008(\bench_v[5] [25]),
        .g1015(\bench_vout[5] [8]),
        .g1016(\bench_v[5] [26]),
        .g1017(\bench_vout[5] [9]),
        .g1080(\bench_v[5] [27]),
        .g1234(\bench_v[5] [28]),
        .g1246(\bench_vout[5] [10]),
        .g1553(\bench_v[5] [29]),
        .g1554(\bench_v[5] [30]),
        .g1724(\bench_vout[5] [11]),
        .g1783(\bench_vout[5] [12]),
        .g1798(\bench_vout[5] [13]),
        .g1804(\bench_vout[5] [14]),
        .g1810(\bench_vout[5] [15]),
        .g1817(\bench_vout[5] [16]),
        .g1824(\bench_vout[5] [17]),
        .g1829(\bench_vout[5] [18]),
        .g1870(\bench_vout[5] [19]),
        .g1871(\bench_vout[5] [20]),
        .g1894(\bench_vout[5] [21]),
        .g1911(\bench_vout[5] [22]),
        .g1944(\bench_vout[5] [23]),
        .g206(\bench_vout[5] [0]),
        .g2662(\bench_vout[5] [24]),
        .g2844(\bench_vout[5] [25]),
        .g2888(\bench_vout[5] [26]),
        .g291(\bench_vout[5] [1]),
        .g3077(\bench_vout[5] [27]),
        .g3096(\bench_vout[5] [28]),
        .g3130(\bench_vout[5] [29]),
        .g3159(\bench_vout[5] [30]),
        .g3191(\bench_vout[5] [31]),
        .g372(\bench_vout[5] [2]),
        .g3829(\bench_vout[5] [32]),
        .g3859(\bench_vout[5] [33]),
        .g3860(\bench_vout[5] [34]),
        .g4267(\bench_vout[5] [35]),
        .g43(\bench_v[5] [0]),
        .g4316(\bench_vout[5] [36]),
        .g4370(\bench_vout[5] [37]),
        .g4371(\bench_vout[5] [38]),
        .g4372(\bench_vout[5] [39]),
        .g4373(\bench_vout[5] [40]),
        .g453(\bench_vout[5] [3]),
        .g4655(\bench_vout[5] [41]),
        .g4657(\bench_vout[5] [42]),
        .g4660(\bench_vout[5] [43]),
        .g4661(\bench_vout[5] [44]),
        .g4663(\bench_vout[5] [45]),
        .g4664(\bench_vout[5] [46]),
        .g49(\bench_v[5] [1]),
        .g5143(\bench_vout[5] [47]),
        .g5164(\bench_vout[5] [48]),
        .g534(\bench_vout[5] [4]),
        .g5571(\bench_vout[5] [49]),
        .g5669(\bench_vout[5] [50]),
        .g5678(\bench_vout[5] [51]),
        .g5682(\bench_vout[5] [52]),
        .g5684(\bench_vout[5] [53]),
        .g5687(\bench_vout[5] [54]),
        .g5729(\bench_vout[5] [55]),
        .g594(\bench_vout[5] [5]),
        .g6207(\bench_vout[5] [56]),
        .g6212(\bench_vout[5] [57]),
        .g6223(\bench_vout[5] [58]),
        .g6236(\bench_vout[5] [59]),
        .g6269(\bench_vout[5] [60]),
        .g633(\bench_v[5] [2]),
        .g634(\bench_v[5] [3]),
        .g635(\bench_v[5] [4]),
        .g6425(\bench_vout[5] [61]),
        .g645(\bench_v[5] [5]),
        .g647(\bench_v[5] [6]),
        .g648(\bench_v[5] [7]),
        .g6648(\bench_vout[5] [62]),
        .g6653(\bench_vout[5] [63]),
        .g6675(\bench_vout[5] [64]),
        .g6849(\bench_vout[5] [65]),
        .g6850(\bench_vout[5] [66]),
        .g6895(\bench_vout[5] [67]),
        .g690(\bench_v[5] [8]),
        .g6909(\bench_vout[5] [68]),
        .g694(\bench_v[5] [9]),
        .g698(\bench_v[5] [10]),
        .g702(\bench_v[5] [11]),
        .g7048(\bench_vout[5] [69]),
        .g7063(\bench_vout[5] [70]),
        .g7103(\bench_vout[5] [71]),
        .g722(\bench_v[5] [12]),
        .g723(\bench_v[5] [13]),
        .g7283(\bench_vout[5] [72]),
        .g7284(\bench_vout[5] [73]),
        .g7285(\bench_vout[5] [74]),
        .g7286(\bench_vout[5] [75]),
        .g7287(\bench_vout[5] [76]),
        .g7288(\bench_vout[5] [77]),
        .g7289(\bench_vout[5] [78]),
        .g7290(\bench_vout[5] [79]),
        .g7291(\bench_vout[5] [80]),
        .g7292(\bench_vout[5] [81]),
        .g7293(\bench_vout[5] [82]),
        .g7294(\bench_vout[5] [83]),
        .g7295(\bench_vout[5] [84]),
        .g7298(\bench_vout[5] [85]),
        .g7423(\bench_vout[5] [86]),
        .g7424(\bench_vout[5] [87]),
        .g7425(\bench_vout[5] [88]),
        .g7474(\bench_vout[5] [89]),
        .g7504(\bench_vout[5] [90]),
        .g7505(\bench_vout[5] [91]),
        .g7506(\bench_vout[5] [92]),
        .g7507(\bench_vout[5] [93]),
        .g7508(\bench_vout[5] [94]),
        .g751(\bench_v[5] [14]),
        .g7514(\bench_vout[5] [95]),
        .g752(\bench_v[5] [15]),
        .g753(\bench_v[5] [16]),
        .g754(\bench_v[5] [17]),
        .g755(\bench_v[5] [18]),
        .g756(\bench_v[5] [19]),
        .g757(\bench_v[5] [20]),
        .g7729(\bench_vout[5] [96]),
        .g7730(\bench_vout[5] [97]),
        .g7731(\bench_vout[5] [98]),
        .g7732(\bench_vout[5] [99]),
        .g781(\bench_v[5] [21]),
        .g785(\bench_vout[5] [6]),
        .g8216(\bench_vout[5] [100]),
        .g8217(\bench_vout[5] [101]),
        .g8218(\bench_vout[5] [102]),
        .g8219(\bench_vout[5] [103]),
        .g8234(\bench_vout[5] [104]),
        .g8661(\bench_vout[5] [105]),
        .g8663(\bench_vout[5] [106]),
        .g8872(\bench_vout[5] [107]),
        .g8958(\bench_vout[5] [108]),
        .g9128(\bench_vout[5] [109]),
        .g9132(\bench_vout[5] [110]),
        .g9204(\bench_vout[5] [111]),
        .g9280(\bench_vout[5] [112]),
        .g9297(\bench_vout[5] [113]),
        .g9299(\bench_vout[5] [114]),
        .g9305(\bench_vout[5] [115]),
        .g9308(\bench_vout[5] [116]),
        .g9310(\bench_vout[5] [117]),
        .g9312(\bench_vout[5] [118]),
        .g9314(\bench_vout[5] [119]),
        .g9378(\bench_vout[5] [120]),
        .g941(\bench_v[5] [22]),
        .g962(\bench_v[5] [23]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][0] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [0]),
        .Q(\bench_vout_reg[6] [0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][100] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [100]),
        .Q(\bench_vout_reg[6] [100]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][101] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [101]),
        .Q(\bench_vout_reg[6] [101]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][102] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [102]),
        .Q(\bench_vout_reg[6] [102]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][103] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [103]),
        .Q(\bench_vout_reg[6] [103]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][104] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [104]),
        .Q(\bench_vout_reg[6] [104]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][105] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [105]),
        .Q(\bench_vout_reg[6] [105]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][106] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [106]),
        .Q(\bench_vout_reg[6] [106]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][107] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [107]),
        .Q(\bench_vout_reg[6] [107]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][108] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [108]),
        .Q(\bench_vout_reg[6] [108]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][109] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [109]),
        .Q(\bench_vout_reg[6] [109]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][10] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [10]),
        .Q(\bench_vout_reg[6] [10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][110] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [110]),
        .Q(\bench_vout_reg[6] [110]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][111] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [111]),
        .Q(\bench_vout_reg[6] [111]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][112] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [112]),
        .Q(\bench_vout_reg[6] [112]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][113] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [113]),
        .Q(\bench_vout_reg[6] [113]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][114] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [114]),
        .Q(\bench_vout_reg[6] [114]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][115] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [115]),
        .Q(\bench_vout_reg[6] [115]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][116] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [116]),
        .Q(\bench_vout_reg[6] [116]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][117] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [117]),
        .Q(\bench_vout_reg[6] [117]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][118] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [118]),
        .Q(\bench_vout_reg[6] [118]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][119] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [119]),
        .Q(\bench_vout_reg[6] [119]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][11] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [11]),
        .Q(\bench_vout_reg[6] [11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][120] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [120]),
        .Q(\bench_vout_reg[6] [120]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][12] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [12]),
        .Q(\bench_vout_reg[6] [12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][13] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [13]),
        .Q(\bench_vout_reg[6] [13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][14] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [14]),
        .Q(\bench_vout_reg[6] [14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][15] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [15]),
        .Q(\bench_vout_reg[6] [15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][16] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [16]),
        .Q(\bench_vout_reg[6] [16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][17] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [17]),
        .Q(\bench_vout_reg[6] [17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][18] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [18]),
        .Q(\bench_vout_reg[6] [18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][19] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [19]),
        .Q(\bench_vout_reg[6] [19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][1] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [1]),
        .Q(\bench_vout_reg[6] [1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][20] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [20]),
        .Q(\bench_vout_reg[6] [20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][21] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [21]),
        .Q(\bench_vout_reg[6] [21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][22] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [22]),
        .Q(\bench_vout_reg[6] [22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][23] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [23]),
        .Q(\bench_vout_reg[6] [23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][24] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [24]),
        .Q(\bench_vout_reg[6] [24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][25] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [25]),
        .Q(\bench_vout_reg[6] [25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][26] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [26]),
        .Q(\bench_vout_reg[6] [26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][27] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [27]),
        .Q(\bench_vout_reg[6] [27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][28] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [28]),
        .Q(\bench_vout_reg[6] [28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][29] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [29]),
        .Q(\bench_vout_reg[6] [29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][2] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [2]),
        .Q(\bench_vout_reg[6] [2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][30] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [30]),
        .Q(\bench_vout_reg[6] [30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][31] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [31]),
        .Q(\bench_vout_reg[6] [31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][32] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [32]),
        .Q(\bench_vout_reg[6] [32]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][33] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [33]),
        .Q(\bench_vout_reg[6] [33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][34] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [34]),
        .Q(\bench_vout_reg[6] [34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][35] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [35]),
        .Q(\bench_vout_reg[6] [35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][36] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [36]),
        .Q(\bench_vout_reg[6] [36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][37] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [37]),
        .Q(\bench_vout_reg[6] [37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][38] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [38]),
        .Q(\bench_vout_reg[6] [38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][39] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [39]),
        .Q(\bench_vout_reg[6] [39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][3] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [3]),
        .Q(\bench_vout_reg[6] [3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][40] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [40]),
        .Q(\bench_vout_reg[6] [40]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][41] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [41]),
        .Q(\bench_vout_reg[6] [41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][42] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [42]),
        .Q(\bench_vout_reg[6] [42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][43] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [43]),
        .Q(\bench_vout_reg[6] [43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][44] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [44]),
        .Q(\bench_vout_reg[6] [44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][45] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [45]),
        .Q(\bench_vout_reg[6] [45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][46] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [46]),
        .Q(\bench_vout_reg[6] [46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][47] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [47]),
        .Q(\bench_vout_reg[6] [47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][48] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [48]),
        .Q(\bench_vout_reg[6] [48]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][49] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [49]),
        .Q(\bench_vout_reg[6] [49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][4] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [4]),
        .Q(\bench_vout_reg[6] [4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][50] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [50]),
        .Q(\bench_vout_reg[6] [50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][51] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [51]),
        .Q(\bench_vout_reg[6] [51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][52] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [52]),
        .Q(\bench_vout_reg[6] [52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][53] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [53]),
        .Q(\bench_vout_reg[6] [53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][54] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [54]),
        .Q(\bench_vout_reg[6] [54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][55] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [55]),
        .Q(\bench_vout_reg[6] [55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][56] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [56]),
        .Q(\bench_vout_reg[6] [56]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][57] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [57]),
        .Q(\bench_vout_reg[6] [57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][58] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [58]),
        .Q(\bench_vout_reg[6] [58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][59] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [59]),
        .Q(\bench_vout_reg[6] [59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][5] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [5]),
        .Q(\bench_vout_reg[6] [5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][60] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [60]),
        .Q(\bench_vout_reg[6] [60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][61] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [61]),
        .Q(\bench_vout_reg[6] [61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][62] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [62]),
        .Q(\bench_vout_reg[6] [62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][63] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [63]),
        .Q(\bench_vout_reg[6] [63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][64] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [64]),
        .Q(\bench_vout_reg[6] [64]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][65] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [65]),
        .Q(\bench_vout_reg[6] [65]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][66] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [66]),
        .Q(\bench_vout_reg[6] [66]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][67] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [67]),
        .Q(\bench_vout_reg[6] [67]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][68] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [68]),
        .Q(\bench_vout_reg[6] [68]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][69] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [69]),
        .Q(\bench_vout_reg[6] [69]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][6] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [6]),
        .Q(\bench_vout_reg[6] [6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][70] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [70]),
        .Q(\bench_vout_reg[6] [70]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][71] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [71]),
        .Q(\bench_vout_reg[6] [71]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][72] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [72]),
        .Q(\bench_vout_reg[6] [72]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][73] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [73]),
        .Q(\bench_vout_reg[6] [73]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][74] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [74]),
        .Q(\bench_vout_reg[6] [74]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][75] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [75]),
        .Q(\bench_vout_reg[6] [75]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][76] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [76]),
        .Q(\bench_vout_reg[6] [76]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][77] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [77]),
        .Q(\bench_vout_reg[6] [77]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][78] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [78]),
        .Q(\bench_vout_reg[6] [78]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][79] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [79]),
        .Q(\bench_vout_reg[6] [79]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][7] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [7]),
        .Q(\bench_vout_reg[6] [7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][80] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [80]),
        .Q(\bench_vout_reg[6] [80]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][81] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [81]),
        .Q(\bench_vout_reg[6] [81]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][82] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [82]),
        .Q(\bench_vout_reg[6] [82]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][83] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [83]),
        .Q(\bench_vout_reg[6] [83]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][84] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [84]),
        .Q(\bench_vout_reg[6] [84]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][85] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [85]),
        .Q(\bench_vout_reg[6] [85]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][86] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [86]),
        .Q(\bench_vout_reg[6] [86]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][87] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [87]),
        .Q(\bench_vout_reg[6] [87]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][88] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [88]),
        .Q(\bench_vout_reg[6] [88]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][89] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [89]),
        .Q(\bench_vout_reg[6] [89]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][8] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [8]),
        .Q(\bench_vout_reg[6] [8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][90] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [90]),
        .Q(\bench_vout_reg[6] [90]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][91] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [91]),
        .Q(\bench_vout_reg[6] [91]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][92] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [92]),
        .Q(\bench_vout_reg[6] [92]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][93] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [93]),
        .Q(\bench_vout_reg[6] [93]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][94] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [94]),
        .Q(\bench_vout_reg[6] [94]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][95] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [95]),
        .Q(\bench_vout_reg[6] [95]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][96] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [96]),
        .Q(\bench_vout_reg[6] [96]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][97] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [97]),
        .Q(\bench_vout_reg[6] [97]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][98] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [98]),
        .Q(\bench_vout_reg[6] [98]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][99] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [99]),
        .Q(\bench_vout_reg[6] [99]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  (* s = "true" *) 
  FDRE #(
    .INIT(1'b0)) 
    \noise_circ_replica[6].bench_vout_reg_reg[6][9] 
       (.C(sysclk),
        .CE(1'b1),
        .D(\bench_vout[6] [9]),
        .Q(\bench_vout_reg[6] [9]),
        .R(1'b0));
  (* KEEP = "true" *) 
  switch_elements_rng \noise_circ_replica[6].lfsr_inst 
       (.clk(sysclk),
        .loadseed_i(loadseed_s),
        .number_o(\random_data_s[6] ),
        .reset(noise_enable_s),
        .seed_i(\seed_s[6] ));
  (* KEEP = "true" *) 
  switch_elements_s13207_bench \noise_circ_replica[6].s13207_bench_inst 
       (.blif_clk_net(sysclk),
        .blif_reset_net(n_noise_enable_s),
        .g1000(\bench_v[6] [24]),
        .g1006(\bench_vout[6] [7]),
        .g1008(\bench_v[6] [25]),
        .g1015(\bench_vout[6] [8]),
        .g1016(\bench_v[6] [26]),
        .g1017(\bench_vout[6] [9]),
        .g1080(\bench_v[6] [27]),
        .g1234(\bench_v[6] [28]),
        .g1246(\bench_vout[6] [10]),
        .g1553(\bench_v[6] [29]),
        .g1554(\bench_v[6] [30]),
        .g1724(\bench_vout[6] [11]),
        .g1783(\bench_vout[6] [12]),
        .g1798(\bench_vout[6] [13]),
        .g1804(\bench_vout[6] [14]),
        .g1810(\bench_vout[6] [15]),
        .g1817(\bench_vout[6] [16]),
        .g1824(\bench_vout[6] [17]),
        .g1829(\bench_vout[6] [18]),
        .g1870(\bench_vout[6] [19]),
        .g1871(\bench_vout[6] [20]),
        .g1894(\bench_vout[6] [21]),
        .g1911(\bench_vout[6] [22]),
        .g1944(\bench_vout[6] [23]),
        .g206(\bench_vout[6] [0]),
        .g2662(\bench_vout[6] [24]),
        .g2844(\bench_vout[6] [25]),
        .g2888(\bench_vout[6] [26]),
        .g291(\bench_vout[6] [1]),
        .g3077(\bench_vout[6] [27]),
        .g3096(\bench_vout[6] [28]),
        .g3130(\bench_vout[6] [29]),
        .g3159(\bench_vout[6] [30]),
        .g3191(\bench_vout[6] [31]),
        .g372(\bench_vout[6] [2]),
        .g3829(\bench_vout[6] [32]),
        .g3859(\bench_vout[6] [33]),
        .g3860(\bench_vout[6] [34]),
        .g4267(\bench_vout[6] [35]),
        .g43(\bench_v[6] [0]),
        .g4316(\bench_vout[6] [36]),
        .g4370(\bench_vout[6] [37]),
        .g4371(\bench_vout[6] [38]),
        .g4372(\bench_vout[6] [39]),
        .g4373(\bench_vout[6] [40]),
        .g453(\bench_vout[6] [3]),
        .g4655(\bench_vout[6] [41]),
        .g4657(\bench_vout[6] [42]),
        .g4660(\bench_vout[6] [43]),
        .g4661(\bench_vout[6] [44]),
        .g4663(\bench_vout[6] [45]),
        .g4664(\bench_vout[6] [46]),
        .g49(\bench_v[6] [1]),
        .g5143(\bench_vout[6] [47]),
        .g5164(\bench_vout[6] [48]),
        .g534(\bench_vout[6] [4]),
        .g5571(\bench_vout[6] [49]),
        .g5669(\bench_vout[6] [50]),
        .g5678(\bench_vout[6] [51]),
        .g5682(\bench_vout[6] [52]),
        .g5684(\bench_vout[6] [53]),
        .g5687(\bench_vout[6] [54]),
        .g5729(\bench_vout[6] [55]),
        .g594(\bench_vout[6] [5]),
        .g6207(\bench_vout[6] [56]),
        .g6212(\bench_vout[6] [57]),
        .g6223(\bench_vout[6] [58]),
        .g6236(\bench_vout[6] [59]),
        .g6269(\bench_vout[6] [60]),
        .g633(\bench_v[6] [2]),
        .g634(\bench_v[6] [3]),
        .g635(\bench_v[6] [4]),
        .g6425(\bench_vout[6] [61]),
        .g645(\bench_v[6] [5]),
        .g647(\bench_v[6] [6]),
        .g648(\bench_v[6] [7]),
        .g6648(\bench_vout[6] [62]),
        .g6653(\bench_vout[6] [63]),
        .g6675(\bench_vout[6] [64]),
        .g6849(\bench_vout[6] [65]),
        .g6850(\bench_vout[6] [66]),
        .g6895(\bench_vout[6] [67]),
        .g690(\bench_v[6] [8]),
        .g6909(\bench_vout[6] [68]),
        .g694(\bench_v[6] [9]),
        .g698(\bench_v[6] [10]),
        .g702(\bench_v[6] [11]),
        .g7048(\bench_vout[6] [69]),
        .g7063(\bench_vout[6] [70]),
        .g7103(\bench_vout[6] [71]),
        .g722(\bench_v[6] [12]),
        .g723(\bench_v[6] [13]),
        .g7283(\bench_vout[6] [72]),
        .g7284(\bench_vout[6] [73]),
        .g7285(\bench_vout[6] [74]),
        .g7286(\bench_vout[6] [75]),
        .g7287(\bench_vout[6] [76]),
        .g7288(\bench_vout[6] [77]),
        .g7289(\bench_vout[6] [78]),
        .g7290(\bench_vout[6] [79]),
        .g7291(\bench_vout[6] [80]),
        .g7292(\bench_vout[6] [81]),
        .g7293(\bench_vout[6] [82]),
        .g7294(\bench_vout[6] [83]),
        .g7295(\bench_vout[6] [84]),
        .g7298(\bench_vout[6] [85]),
        .g7423(\bench_vout[6] [86]),
        .g7424(\bench_vout[6] [87]),
        .g7425(\bench_vout[6] [88]),
        .g7474(\bench_vout[6] [89]),
        .g7504(\bench_vout[6] [90]),
        .g7505(\bench_vout[6] [91]),
        .g7506(\bench_vout[6] [92]),
        .g7507(\bench_vout[6] [93]),
        .g7508(\bench_vout[6] [94]),
        .g751(\bench_v[6] [14]),
        .g7514(\bench_vout[6] [95]),
        .g752(\bench_v[6] [15]),
        .g753(\bench_v[6] [16]),
        .g754(\bench_v[6] [17]),
        .g755(\bench_v[6] [18]),
        .g756(\bench_v[6] [19]),
        .g757(\bench_v[6] [20]),
        .g7729(\bench_vout[6] [96]),
        .g7730(\bench_vout[6] [97]),
        .g7731(\bench_vout[6] [98]),
        .g7732(\bench_vout[6] [99]),
        .g781(\bench_v[6] [21]),
        .g785(\bench_vout[6] [6]),
        .g8216(\bench_vout[6] [100]),
        .g8217(\bench_vout[6] [101]),
        .g8218(\bench_vout[6] [102]),
        .g8219(\bench_vout[6] [103]),
        .g8234(\bench_vout[6] [104]),
        .g8661(\bench_vout[6] [105]),
        .g8663(\bench_vout[6] [106]),
        .g8872(\bench_vout[6] [107]),
        .g8958(\bench_vout[6] [108]),
        .g9128(\bench_vout[6] [109]),
        .g9132(\bench_vout[6] [110]),
        .g9204(\bench_vout[6] [111]),
        .g9280(\bench_vout[6] [112]),
        .g9297(\bench_vout[6] [113]),
        .g9299(\bench_vout[6] [114]),
        .g9305(\bench_vout[6] [115]),
        .g9308(\bench_vout[6] [116]),
        .g9310(\bench_vout[6] [117]),
        .g9312(\bench_vout[6] [118]),
        .g9314(\bench_vout[6] [119]),
        .g9378(\bench_vout[6] [120]),
        .g941(\bench_v[6] [22]),
        .g962(\bench_v[6] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst 
       (.I0(\random_data_s[0] [30]),
        .O(\bench_v[0] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__0 
       (.I0(\random_data_s[0] [29]),
        .O(\bench_v[0] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__1 
       (.I0(\random_data_s[0] [28]),
        .O(\bench_v[0] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__10 
       (.I0(\random_data_s[0] [19]),
        .O(\bench_v[0] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__11 
       (.I0(\random_data_s[0] [18]),
        .O(\bench_v[0] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__12 
       (.I0(\random_data_s[0] [17]),
        .O(\bench_v[0] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__13 
       (.I0(\random_data_s[0] [16]),
        .O(\bench_v[0] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__14 
       (.I0(\random_data_s[0] [15]),
        .O(\bench_v[0] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__15 
       (.I0(\random_data_s[0] [14]),
        .O(\bench_v[0] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__16 
       (.I0(\random_data_s[0] [13]),
        .O(\bench_v[0] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__17 
       (.I0(\random_data_s[0] [12]),
        .O(\bench_v[0] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__18 
       (.I0(\random_data_s[0] [11]),
        .O(\bench_v[0] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__19 
       (.I0(\random_data_s[0] [10]),
        .O(\bench_v[0] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__2 
       (.I0(\random_data_s[0] [27]),
        .O(\bench_v[0] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__20 
       (.I0(\random_data_s[0] [9]),
        .O(\bench_v[0] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__21 
       (.I0(\random_data_s[0] [8]),
        .O(\bench_v[0] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__22 
       (.I0(\random_data_s[0] [7]),
        .O(\bench_v[0] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__23 
       (.I0(\random_data_s[0] [6]),
        .O(\bench_v[0] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__24 
       (.I0(\random_data_s[0] [5]),
        .O(\bench_v[0] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__25 
       (.I0(\random_data_s[0] [4]),
        .O(\bench_v[0] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__26 
       (.I0(\random_data_s[0] [3]),
        .O(\bench_v[0] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__27 
       (.I0(\random_data_s[0] [2]),
        .O(\bench_v[0] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__28 
       (.I0(\random_data_s[0] [1]),
        .O(\bench_v[0] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__29 
       (.I0(\random_data_s[0] [0]),
        .O(\bench_v[0] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__3 
       (.I0(\random_data_s[0] [26]),
        .O(\bench_v[0] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__4 
       (.I0(\random_data_s[0] [25]),
        .O(\bench_v[0] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__5 
       (.I0(\random_data_s[0] [24]),
        .O(\bench_v[0] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__6 
       (.I0(\random_data_s[0] [23]),
        .O(\bench_v[0] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__7 
       (.I0(\random_data_s[0] [22]),
        .O(\bench_v[0] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__8 
       (.I0(\random_data_s[0] [21]),
        .O(\bench_v[0] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[0]_inst__9 
       (.I0(\random_data_s[0] [20]),
        .O(\bench_v[0] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst 
       (.I0(\random_data_s[1] [30]),
        .O(\bench_v[1] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__0 
       (.I0(\random_data_s[1] [29]),
        .O(\bench_v[1] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__1 
       (.I0(\random_data_s[1] [28]),
        .O(\bench_v[1] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__10 
       (.I0(\random_data_s[1] [19]),
        .O(\bench_v[1] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__11 
       (.I0(\random_data_s[1] [18]),
        .O(\bench_v[1] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__12 
       (.I0(\random_data_s[1] [17]),
        .O(\bench_v[1] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__13 
       (.I0(\random_data_s[1] [16]),
        .O(\bench_v[1] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__14 
       (.I0(\random_data_s[1] [15]),
        .O(\bench_v[1] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__15 
       (.I0(\random_data_s[1] [14]),
        .O(\bench_v[1] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__16 
       (.I0(\random_data_s[1] [13]),
        .O(\bench_v[1] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__17 
       (.I0(\random_data_s[1] [12]),
        .O(\bench_v[1] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__18 
       (.I0(\random_data_s[1] [11]),
        .O(\bench_v[1] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__19 
       (.I0(\random_data_s[1] [10]),
        .O(\bench_v[1] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__2 
       (.I0(\random_data_s[1] [27]),
        .O(\bench_v[1] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__20 
       (.I0(\random_data_s[1] [9]),
        .O(\bench_v[1] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__21 
       (.I0(\random_data_s[1] [8]),
        .O(\bench_v[1] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__22 
       (.I0(\random_data_s[1] [7]),
        .O(\bench_v[1] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__23 
       (.I0(\random_data_s[1] [6]),
        .O(\bench_v[1] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__24 
       (.I0(\random_data_s[1] [5]),
        .O(\bench_v[1] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__25 
       (.I0(\random_data_s[1] [4]),
        .O(\bench_v[1] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__26 
       (.I0(\random_data_s[1] [3]),
        .O(\bench_v[1] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__27 
       (.I0(\random_data_s[1] [2]),
        .O(\bench_v[1] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__28 
       (.I0(\random_data_s[1] [1]),
        .O(\bench_v[1] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__29 
       (.I0(\random_data_s[1] [0]),
        .O(\bench_v[1] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__3 
       (.I0(\random_data_s[1] [26]),
        .O(\bench_v[1] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__4 
       (.I0(\random_data_s[1] [25]),
        .O(\bench_v[1] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__5 
       (.I0(\random_data_s[1] [24]),
        .O(\bench_v[1] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__6 
       (.I0(\random_data_s[1] [23]),
        .O(\bench_v[1] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__7 
       (.I0(\random_data_s[1] [22]),
        .O(\bench_v[1] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__8 
       (.I0(\random_data_s[1] [21]),
        .O(\bench_v[1] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[1]_inst__9 
       (.I0(\random_data_s[1] [20]),
        .O(\bench_v[1] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst 
       (.I0(\random_data_s[2] [30]),
        .O(\bench_v[2] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__0 
       (.I0(\random_data_s[2] [29]),
        .O(\bench_v[2] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__1 
       (.I0(\random_data_s[2] [28]),
        .O(\bench_v[2] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__10 
       (.I0(\random_data_s[2] [19]),
        .O(\bench_v[2] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__11 
       (.I0(\random_data_s[2] [18]),
        .O(\bench_v[2] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__12 
       (.I0(\random_data_s[2] [17]),
        .O(\bench_v[2] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__13 
       (.I0(\random_data_s[2] [16]),
        .O(\bench_v[2] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__14 
       (.I0(\random_data_s[2] [15]),
        .O(\bench_v[2] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__15 
       (.I0(\random_data_s[2] [14]),
        .O(\bench_v[2] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__16 
       (.I0(\random_data_s[2] [13]),
        .O(\bench_v[2] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__17 
       (.I0(\random_data_s[2] [12]),
        .O(\bench_v[2] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__18 
       (.I0(\random_data_s[2] [11]),
        .O(\bench_v[2] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__19 
       (.I0(\random_data_s[2] [10]),
        .O(\bench_v[2] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__2 
       (.I0(\random_data_s[2] [27]),
        .O(\bench_v[2] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__20 
       (.I0(\random_data_s[2] [9]),
        .O(\bench_v[2] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__21 
       (.I0(\random_data_s[2] [8]),
        .O(\bench_v[2] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__22 
       (.I0(\random_data_s[2] [7]),
        .O(\bench_v[2] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__23 
       (.I0(\random_data_s[2] [6]),
        .O(\bench_v[2] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__24 
       (.I0(\random_data_s[2] [5]),
        .O(\bench_v[2] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__25 
       (.I0(\random_data_s[2] [4]),
        .O(\bench_v[2] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__26 
       (.I0(\random_data_s[2] [3]),
        .O(\bench_v[2] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__27 
       (.I0(\random_data_s[2] [2]),
        .O(\bench_v[2] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__28 
       (.I0(\random_data_s[2] [1]),
        .O(\bench_v[2] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__29 
       (.I0(\random_data_s[2] [0]),
        .O(\bench_v[2] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__3 
       (.I0(\random_data_s[2] [26]),
        .O(\bench_v[2] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__4 
       (.I0(\random_data_s[2] [25]),
        .O(\bench_v[2] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__5 
       (.I0(\random_data_s[2] [24]),
        .O(\bench_v[2] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__6 
       (.I0(\random_data_s[2] [23]),
        .O(\bench_v[2] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__7 
       (.I0(\random_data_s[2] [22]),
        .O(\bench_v[2] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__8 
       (.I0(\random_data_s[2] [21]),
        .O(\bench_v[2] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[2]_inst__9 
       (.I0(\random_data_s[2] [20]),
        .O(\bench_v[2] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst 
       (.I0(\random_data_s[3] [30]),
        .O(\bench_v[3] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__0 
       (.I0(\random_data_s[3] [29]),
        .O(\bench_v[3] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__1 
       (.I0(\random_data_s[3] [28]),
        .O(\bench_v[3] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__10 
       (.I0(\random_data_s[3] [19]),
        .O(\bench_v[3] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__11 
       (.I0(\random_data_s[3] [18]),
        .O(\bench_v[3] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__12 
       (.I0(\random_data_s[3] [17]),
        .O(\bench_v[3] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__13 
       (.I0(\random_data_s[3] [16]),
        .O(\bench_v[3] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__14 
       (.I0(\random_data_s[3] [15]),
        .O(\bench_v[3] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__15 
       (.I0(\random_data_s[3] [14]),
        .O(\bench_v[3] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__16 
       (.I0(\random_data_s[3] [13]),
        .O(\bench_v[3] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__17 
       (.I0(\random_data_s[3] [12]),
        .O(\bench_v[3] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__18 
       (.I0(\random_data_s[3] [11]),
        .O(\bench_v[3] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__19 
       (.I0(\random_data_s[3] [10]),
        .O(\bench_v[3] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__2 
       (.I0(\random_data_s[3] [27]),
        .O(\bench_v[3] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__20 
       (.I0(\random_data_s[3] [9]),
        .O(\bench_v[3] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__21 
       (.I0(\random_data_s[3] [8]),
        .O(\bench_v[3] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__22 
       (.I0(\random_data_s[3] [7]),
        .O(\bench_v[3] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__23 
       (.I0(\random_data_s[3] [6]),
        .O(\bench_v[3] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__24 
       (.I0(\random_data_s[3] [5]),
        .O(\bench_v[3] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__25 
       (.I0(\random_data_s[3] [4]),
        .O(\bench_v[3] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__26 
       (.I0(\random_data_s[3] [3]),
        .O(\bench_v[3] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__27 
       (.I0(\random_data_s[3] [2]),
        .O(\bench_v[3] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__28 
       (.I0(\random_data_s[3] [1]),
        .O(\bench_v[3] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__29 
       (.I0(\random_data_s[3] [0]),
        .O(\bench_v[3] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__3 
       (.I0(\random_data_s[3] [26]),
        .O(\bench_v[3] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__4 
       (.I0(\random_data_s[3] [25]),
        .O(\bench_v[3] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__5 
       (.I0(\random_data_s[3] [24]),
        .O(\bench_v[3] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__6 
       (.I0(\random_data_s[3] [23]),
        .O(\bench_v[3] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__7 
       (.I0(\random_data_s[3] [22]),
        .O(\bench_v[3] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__8 
       (.I0(\random_data_s[3] [21]),
        .O(\bench_v[3] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[3]_inst__9 
       (.I0(\random_data_s[3] [20]),
        .O(\bench_v[3] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst 
       (.I0(\random_data_s[4] [30]),
        .O(\bench_v[4] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__0 
       (.I0(\random_data_s[4] [29]),
        .O(\bench_v[4] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__1 
       (.I0(\random_data_s[4] [28]),
        .O(\bench_v[4] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__10 
       (.I0(\random_data_s[4] [19]),
        .O(\bench_v[4] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__11 
       (.I0(\random_data_s[4] [18]),
        .O(\bench_v[4] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__12 
       (.I0(\random_data_s[4] [17]),
        .O(\bench_v[4] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__13 
       (.I0(\random_data_s[4] [16]),
        .O(\bench_v[4] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__14 
       (.I0(\random_data_s[4] [15]),
        .O(\bench_v[4] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__15 
       (.I0(\random_data_s[4] [14]),
        .O(\bench_v[4] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__16 
       (.I0(\random_data_s[4] [13]),
        .O(\bench_v[4] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__17 
       (.I0(\random_data_s[4] [12]),
        .O(\bench_v[4] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__18 
       (.I0(\random_data_s[4] [11]),
        .O(\bench_v[4] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__19 
       (.I0(\random_data_s[4] [10]),
        .O(\bench_v[4] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__2 
       (.I0(\random_data_s[4] [27]),
        .O(\bench_v[4] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__20 
       (.I0(\random_data_s[4] [9]),
        .O(\bench_v[4] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__21 
       (.I0(\random_data_s[4] [8]),
        .O(\bench_v[4] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__22 
       (.I0(\random_data_s[4] [7]),
        .O(\bench_v[4] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__23 
       (.I0(\random_data_s[4] [6]),
        .O(\bench_v[4] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__24 
       (.I0(\random_data_s[4] [5]),
        .O(\bench_v[4] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__25 
       (.I0(\random_data_s[4] [4]),
        .O(\bench_v[4] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__26 
       (.I0(\random_data_s[4] [3]),
        .O(\bench_v[4] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__27 
       (.I0(\random_data_s[4] [2]),
        .O(\bench_v[4] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__28 
       (.I0(\random_data_s[4] [1]),
        .O(\bench_v[4] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__29 
       (.I0(\random_data_s[4] [0]),
        .O(\bench_v[4] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__3 
       (.I0(\random_data_s[4] [26]),
        .O(\bench_v[4] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__4 
       (.I0(\random_data_s[4] [25]),
        .O(\bench_v[4] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__5 
       (.I0(\random_data_s[4] [24]),
        .O(\bench_v[4] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__6 
       (.I0(\random_data_s[4] [23]),
        .O(\bench_v[4] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__7 
       (.I0(\random_data_s[4] [22]),
        .O(\bench_v[4] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__8 
       (.I0(\random_data_s[4] [21]),
        .O(\bench_v[4] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[4]_inst__9 
       (.I0(\random_data_s[4] [20]),
        .O(\bench_v[4] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst 
       (.I0(\random_data_s[5] [30]),
        .O(\bench_v[5] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__0 
       (.I0(\random_data_s[5] [29]),
        .O(\bench_v[5] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__1 
       (.I0(\random_data_s[5] [28]),
        .O(\bench_v[5] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__10 
       (.I0(\random_data_s[5] [19]),
        .O(\bench_v[5] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__11 
       (.I0(\random_data_s[5] [18]),
        .O(\bench_v[5] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__12 
       (.I0(\random_data_s[5] [17]),
        .O(\bench_v[5] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__13 
       (.I0(\random_data_s[5] [16]),
        .O(\bench_v[5] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__14 
       (.I0(\random_data_s[5] [15]),
        .O(\bench_v[5] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__15 
       (.I0(\random_data_s[5] [14]),
        .O(\bench_v[5] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__16 
       (.I0(\random_data_s[5] [13]),
        .O(\bench_v[5] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__17 
       (.I0(\random_data_s[5] [12]),
        .O(\bench_v[5] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__18 
       (.I0(\random_data_s[5] [11]),
        .O(\bench_v[5] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__19 
       (.I0(\random_data_s[5] [10]),
        .O(\bench_v[5] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__2 
       (.I0(\random_data_s[5] [27]),
        .O(\bench_v[5] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__20 
       (.I0(\random_data_s[5] [9]),
        .O(\bench_v[5] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__21 
       (.I0(\random_data_s[5] [8]),
        .O(\bench_v[5] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__22 
       (.I0(\random_data_s[5] [7]),
        .O(\bench_v[5] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__23 
       (.I0(\random_data_s[5] [6]),
        .O(\bench_v[5] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__24 
       (.I0(\random_data_s[5] [5]),
        .O(\bench_v[5] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__25 
       (.I0(\random_data_s[5] [4]),
        .O(\bench_v[5] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__26 
       (.I0(\random_data_s[5] [3]),
        .O(\bench_v[5] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__27 
       (.I0(\random_data_s[5] [2]),
        .O(\bench_v[5] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__28 
       (.I0(\random_data_s[5] [1]),
        .O(\bench_v[5] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__29 
       (.I0(\random_data_s[5] [0]),
        .O(\bench_v[5] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__3 
       (.I0(\random_data_s[5] [26]),
        .O(\bench_v[5] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__4 
       (.I0(\random_data_s[5] [25]),
        .O(\bench_v[5] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__5 
       (.I0(\random_data_s[5] [24]),
        .O(\bench_v[5] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__6 
       (.I0(\random_data_s[5] [23]),
        .O(\bench_v[5] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__7 
       (.I0(\random_data_s[5] [22]),
        .O(\bench_v[5] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__8 
       (.I0(\random_data_s[5] [21]),
        .O(\bench_v[5] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[5]_inst__9 
       (.I0(\random_data_s[5] [20]),
        .O(\bench_v[5] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst 
       (.I0(\random_data_s[6] [30]),
        .O(\bench_v[6] [30]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__0 
       (.I0(\random_data_s[6] [29]),
        .O(\bench_v[6] [29]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__1 
       (.I0(\random_data_s[6] [28]),
        .O(\bench_v[6] [28]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__10 
       (.I0(\random_data_s[6] [19]),
        .O(\bench_v[6] [19]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__11 
       (.I0(\random_data_s[6] [18]),
        .O(\bench_v[6] [18]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__12 
       (.I0(\random_data_s[6] [17]),
        .O(\bench_v[6] [17]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__13 
       (.I0(\random_data_s[6] [16]),
        .O(\bench_v[6] [16]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__14 
       (.I0(\random_data_s[6] [15]),
        .O(\bench_v[6] [15]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__15 
       (.I0(\random_data_s[6] [14]),
        .O(\bench_v[6] [14]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__16 
       (.I0(\random_data_s[6] [13]),
        .O(\bench_v[6] [13]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__17 
       (.I0(\random_data_s[6] [12]),
        .O(\bench_v[6] [12]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__18 
       (.I0(\random_data_s[6] [11]),
        .O(\bench_v[6] [11]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__19 
       (.I0(\random_data_s[6] [10]),
        .O(\bench_v[6] [10]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__2 
       (.I0(\random_data_s[6] [27]),
        .O(\bench_v[6] [27]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__20 
       (.I0(\random_data_s[6] [9]),
        .O(\bench_v[6] [9]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__21 
       (.I0(\random_data_s[6] [8]),
        .O(\bench_v[6] [8]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__22 
       (.I0(\random_data_s[6] [7]),
        .O(\bench_v[6] [7]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__23 
       (.I0(\random_data_s[6] [6]),
        .O(\bench_v[6] [6]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__24 
       (.I0(\random_data_s[6] [5]),
        .O(\bench_v[6] [5]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__25 
       (.I0(\random_data_s[6] [4]),
        .O(\bench_v[6] [4]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__26 
       (.I0(\random_data_s[6] [3]),
        .O(\bench_v[6] [3]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__27 
       (.I0(\random_data_s[6] [2]),
        .O(\bench_v[6] [2]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__28 
       (.I0(\random_data_s[6] [1]),
        .O(\bench_v[6] [1]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__29 
       (.I0(\random_data_s[6] [0]),
        .O(\bench_v[6] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__3 
       (.I0(\random_data_s[6] [26]),
        .O(\bench_v[6] [26]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__4 
       (.I0(\random_data_s[6] [25]),
        .O(\bench_v[6] [25]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__5 
       (.I0(\random_data_s[6] [24]),
        .O(\bench_v[6] [24]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__6 
       (.I0(\random_data_s[6] [23]),
        .O(\bench_v[6] [23]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__7 
       (.I0(\random_data_s[6] [22]),
        .O(\bench_v[6] [22]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__8 
       (.I0(\random_data_s[6] [21]),
        .O(\bench_v[6] [21]));
  LUT1 #(
    .INIT(2'h2)) 
    \random_data_s[6]_inst__9 
       (.I0(\random_data_s[6] [20]),
        .O(\bench_v[6] [20]));
  LUT1 #(
    .INIT(2'h2)) 
    \seed_s[0]_inst 
       (.I0(\seed_s[6] [0]),
        .O(\seed_s[0] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \seed_s[1]_inst 
       (.I0(\seed_s[6] [0]),
        .O(\seed_s[1] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \seed_s[2]_inst 
       (.I0(\seed_s[6] [0]),
        .O(\seed_s[2] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \seed_s[3]_inst 
       (.I0(\seed_s[6] [0]),
        .O(\seed_s[3] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \seed_s[4]_inst 
       (.I0(\seed_s[6] [0]),
        .O(\seed_s[4] [0]));
  LUT1 #(
    .INIT(2'h2)) 
    \seed_s[5]_inst 
       (.I0(\seed_s[6] [0]),
        .O(\seed_s[5] [0]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng__1
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng__2
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng__3
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng__4
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng__5
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "rng" *) 
module switch_elements_rng__6
   (clk,
    reset,
    loadseed_i,
    seed_i,
    number_o);
  input clk;
  input reset;
  input loadseed_i;
  input [31:0]seed_i;
  output [31:0]number_o;

  wire \CASR_reg_reg_n_0_[0] ;
  wire \LFSR_reg[0]_i_1_n_0 ;
  wire \LFSR_reg[10]_i_1_n_0 ;
  wire \LFSR_reg[11]_i_1_n_0 ;
  wire \LFSR_reg[12]_i_1_n_0 ;
  wire \LFSR_reg[13]_i_1_n_0 ;
  wire \LFSR_reg[14]_i_1_n_0 ;
  wire \LFSR_reg[15]_i_1_n_0 ;
  wire \LFSR_reg[16]_i_1_n_0 ;
  wire \LFSR_reg[17]_i_1_n_0 ;
  wire \LFSR_reg[18]_i_1_n_0 ;
  wire \LFSR_reg[19]_i_1_n_0 ;
  wire \LFSR_reg[1]_i_1_n_0 ;
  wire \LFSR_reg[20]_i_1_n_0 ;
  wire \LFSR_reg[21]_i_1_n_0 ;
  wire \LFSR_reg[22]_i_1_n_0 ;
  wire \LFSR_reg[23]_i_1_n_0 ;
  wire \LFSR_reg[24]_i_1_n_0 ;
  wire \LFSR_reg[25]_i_1_n_0 ;
  wire \LFSR_reg[26]_i_1_n_0 ;
  wire \LFSR_reg[27]_i_1_n_0 ;
  wire \LFSR_reg[28]_i_1_n_0 ;
  wire \LFSR_reg[29]_i_1_n_0 ;
  wire \LFSR_reg[2]_i_1_n_0 ;
  wire \LFSR_reg[30]_i_1_n_0 ;
  wire \LFSR_reg[31]_i_1_n_0 ;
  wire \LFSR_reg[32]_i_1_n_0 ;
  wire \LFSR_reg[33]_i_1_n_0 ;
  wire \LFSR_reg[34]_i_1_n_0 ;
  wire \LFSR_reg[35]_i_1_n_0 ;
  wire \LFSR_reg[36]_i_1_n_0 ;
  wire \LFSR_reg[37]_i_1_n_0 ;
  wire \LFSR_reg[38]_i_1_n_0 ;
  wire \LFSR_reg[39]_i_1_n_0 ;
  wire \LFSR_reg[3]_i_1_n_0 ;
  wire \LFSR_reg[40]_i_1_n_0 ;
  wire \LFSR_reg[41]_i_1_n_0 ;
  wire \LFSR_reg[42]_i_1_n_0 ;
  wire \LFSR_reg[4]_i_1_n_0 ;
  wire \LFSR_reg[5]_i_1_n_0 ;
  wire \LFSR_reg[6]_i_1_n_0 ;
  wire \LFSR_reg[7]_i_1_n_0 ;
  wire \LFSR_reg[8]_i_1_n_0 ;
  wire \LFSR_reg[9]_i_1_n_0 ;
  wire \LFSR_reg_reg_n_0_[0] ;
  wire \LFSR_reg_reg_n_0_[10] ;
  wire \LFSR_reg_reg_n_0_[11] ;
  wire \LFSR_reg_reg_n_0_[12] ;
  wire \LFSR_reg_reg_n_0_[13] ;
  wire \LFSR_reg_reg_n_0_[14] ;
  wire \LFSR_reg_reg_n_0_[15] ;
  wire \LFSR_reg_reg_n_0_[16] ;
  wire \LFSR_reg_reg_n_0_[17] ;
  wire \LFSR_reg_reg_n_0_[18] ;
  wire \LFSR_reg_reg_n_0_[1] ;
  wire \LFSR_reg_reg_n_0_[20] ;
  wire \LFSR_reg_reg_n_0_[21] ;
  wire \LFSR_reg_reg_n_0_[22] ;
  wire \LFSR_reg_reg_n_0_[23] ;
  wire \LFSR_reg_reg_n_0_[24] ;
  wire \LFSR_reg_reg_n_0_[25] ;
  wire \LFSR_reg_reg_n_0_[26] ;
  wire \LFSR_reg_reg_n_0_[27] ;
  wire \LFSR_reg_reg_n_0_[28] ;
  wire \LFSR_reg_reg_n_0_[29] ;
  wire \LFSR_reg_reg_n_0_[2] ;
  wire \LFSR_reg_reg_n_0_[30] ;
  wire \LFSR_reg_reg_n_0_[31] ;
  wire \LFSR_reg_reg_n_0_[32] ;
  wire \LFSR_reg_reg_n_0_[33] ;
  wire \LFSR_reg_reg_n_0_[34] ;
  wire \LFSR_reg_reg_n_0_[35] ;
  wire \LFSR_reg_reg_n_0_[36] ;
  wire \LFSR_reg_reg_n_0_[37] ;
  wire \LFSR_reg_reg_n_0_[38] ;
  wire \LFSR_reg_reg_n_0_[39] ;
  wire \LFSR_reg_reg_n_0_[3] ;
  wire \LFSR_reg_reg_n_0_[41] ;
  wire \LFSR_reg_reg_n_0_[4] ;
  wire \LFSR_reg_reg_n_0_[5] ;
  wire \LFSR_reg_reg_n_0_[6] ;
  wire \LFSR_reg_reg_n_0_[7] ;
  wire \LFSR_reg_reg_n_0_[8] ;
  wire \LFSR_reg_reg_n_0_[9] ;
  wire clk;
  wire loadseed_i;
  wire [31:0]number_o;
  wire \number_o[0]_i_1_n_0 ;
  wire \number_o[10]_i_1_n_0 ;
  wire \number_o[11]_i_1_n_0 ;
  wire \number_o[12]_i_1_n_0 ;
  wire \number_o[13]_i_1_n_0 ;
  wire \number_o[14]_i_1_n_0 ;
  wire \number_o[15]_i_1_n_0 ;
  wire \number_o[16]_i_1_n_0 ;
  wire \number_o[17]_i_1_n_0 ;
  wire \number_o[18]_i_1_n_0 ;
  wire \number_o[19]_i_1_n_0 ;
  wire \number_o[1]_i_1_n_0 ;
  wire \number_o[20]_i_1_n_0 ;
  wire \number_o[21]_i_1_n_0 ;
  wire \number_o[22]_i_1_n_0 ;
  wire \number_o[23]_i_1_n_0 ;
  wire \number_o[24]_i_1_n_0 ;
  wire \number_o[25]_i_1_n_0 ;
  wire \number_o[26]_i_1_n_0 ;
  wire \number_o[27]_i_1_n_0 ;
  wire \number_o[28]_i_1_n_0 ;
  wire \number_o[29]_i_1_n_0 ;
  wire \number_o[2]_i_1_n_0 ;
  wire \number_o[30]_i_1_n_0 ;
  wire \number_o[31]_i_1_n_0 ;
  wire \number_o[31]_i_2_n_0 ;
  wire \number_o[3]_i_1_n_0 ;
  wire \number_o[4]_i_1_n_0 ;
  wire \number_o[5]_i_1_n_0 ;
  wire \number_o[6]_i_1_n_0 ;
  wire \number_o[7]_i_1_n_0 ;
  wire \number_o[8]_i_1_n_0 ;
  wire \number_o[9]_i_1_n_0 ;
  wire p_0_in;
  wire p_0_in28_in;
  wire [36:0]p_0_in__0;
  wire p_10_in;
  wire p_11_in;
  wire p_12_in;
  wire p_13_in;
  wire p_14_in;
  wire p_15_in;
  wire p_16_in;
  wire p_17_in;
  wire p_18_in;
  wire p_19_in;
  wire p_1_in;
  wire p_1_in0_in;
  wire p_1_in26_in;
  wire p_20_in;
  wire p_21_in;
  wire p_22_in;
  wire p_23_in;
  wire p_24_in;
  wire p_25_in;
  wire p_26_in;
  wire p_27_in;
  wire p_28_in;
  wire p_29_in;
  wire p_2_in;
  wire p_30_in;
  wire p_31_in;
  wire p_32_in;
  wire p_33_in;
  wire p_34_in;
  wire p_35_in;
  wire p_36_in;
  wire p_3_in;
  wire p_4_in;
  wire p_6_in;
  wire p_7_in;
  wire p_8_in;
  wire p_9_in;
  wire reset;
  wire [31:0]seed_i;

  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(p_2_in),
        .I2(p_3_in),
        .I3(loadseed_i),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(p_14_in),
        .I2(p_12_in),
        .I3(loadseed_i),
        .O(p_0_in__0[10]));
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(p_15_in),
        .I2(p_13_in),
        .I3(loadseed_i),
        .O(p_0_in__0[11]));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(p_16_in),
        .I2(p_14_in),
        .I3(loadseed_i),
        .O(p_0_in__0[12]));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(p_17_in),
        .I2(p_15_in),
        .I3(loadseed_i),
        .O(p_0_in__0[13]));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(p_18_in),
        .I2(p_16_in),
        .I3(loadseed_i),
        .O(p_0_in__0[14]));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(p_19_in),
        .I2(p_17_in),
        .I3(loadseed_i),
        .O(p_0_in__0[15]));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(p_20_in),
        .I2(p_18_in),
        .I3(loadseed_i),
        .O(p_0_in__0[16]));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(p_21_in),
        .I2(p_19_in),
        .I3(loadseed_i),
        .O(p_0_in__0[17]));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(p_22_in),
        .I2(p_20_in),
        .I3(loadseed_i),
        .O(p_0_in__0[18]));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(p_23_in),
        .I2(p_21_in),
        .I3(loadseed_i),
        .O(p_0_in__0[19]));
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(p_4_in),
        .I2(\CASR_reg_reg_n_0_[0] ),
        .I3(loadseed_i),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(p_24_in),
        .I2(p_22_in),
        .I3(loadseed_i),
        .O(p_0_in__0[20]));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(p_25_in),
        .I2(p_23_in),
        .I3(loadseed_i),
        .O(p_0_in__0[21]));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(p_26_in),
        .I2(p_24_in),
        .I3(loadseed_i),
        .O(p_0_in__0[22]));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(p_27_in),
        .I2(p_25_in),
        .I3(loadseed_i),
        .O(p_0_in__0[23]));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(p_28_in),
        .I2(p_26_in),
        .I3(loadseed_i),
        .O(p_0_in__0[24]));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(p_1_in26_in),
        .I2(p_27_in),
        .I3(loadseed_i),
        .O(p_0_in__0[25]));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(p_0_in28_in),
        .I2(p_28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[26]));
  LUT5 #(
    .INIT(32'hAAAAC33C)) 
    \CASR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(p_0_in28_in),
        .I2(p_1_in26_in),
        .I3(p_29_in),
        .I4(loadseed_i),
        .O(p_0_in__0[27]));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(p_30_in),
        .I2(p_0_in28_in),
        .I3(loadseed_i),
        .O(p_0_in__0[28]));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(p_31_in),
        .I2(p_29_in),
        .I3(loadseed_i),
        .O(p_0_in__0[29]));
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(p_6_in),
        .I2(p_2_in),
        .I3(loadseed_i),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(p_32_in),
        .I2(p_30_in),
        .I3(loadseed_i),
        .O(p_0_in__0[30]));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(p_33_in),
        .I2(p_31_in),
        .I3(loadseed_i),
        .O(p_0_in__0[31]));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[32]_i_1 
       (.I0(p_32_in),
        .I1(p_34_in),
        .I2(loadseed_i),
        .O(p_0_in__0[32]));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[33]_i_1 
       (.I0(p_33_in),
        .I1(p_35_in),
        .I2(loadseed_i),
        .O(p_0_in__0[33]));
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[34]_i_1 
       (.I0(p_34_in),
        .I1(p_36_in),
        .I2(loadseed_i),
        .O(p_0_in__0[34]));
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[35]_i_1 
       (.I0(p_35_in),
        .I1(p_3_in),
        .I2(loadseed_i),
        .O(p_0_in__0[35]));
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \CASR_reg[36]_i_1 
       (.I0(p_36_in),
        .I1(\CASR_reg_reg_n_0_[0] ),
        .I2(loadseed_i),
        .O(p_0_in__0[36]));
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(p_7_in),
        .I2(p_4_in),
        .I3(loadseed_i),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(p_8_in),
        .I2(p_6_in),
        .I3(loadseed_i),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(p_9_in),
        .I2(p_7_in),
        .I3(loadseed_i),
        .O(p_0_in__0[5]));
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(p_10_in),
        .I2(p_8_in),
        .I3(loadseed_i),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(p_11_in),
        .I2(p_9_in),
        .I3(loadseed_i),
        .O(p_0_in__0[7]));
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(p_12_in),
        .I2(p_10_in),
        .I3(loadseed_i),
        .O(p_0_in__0[8]));
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT4 #(
    .INIT(16'hAA3C)) 
    \CASR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(p_13_in),
        .I2(p_11_in),
        .I3(loadseed_i),
        .O(p_0_in__0[9]));
  FDPE #(
    .INIT(1'b1)) 
    \CASR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\CASR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[10]),
        .Q(p_13_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[11]),
        .Q(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[12]),
        .Q(p_15_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[13]),
        .Q(p_16_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[14]),
        .Q(p_17_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[15]),
        .Q(p_18_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[16]),
        .Q(p_19_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[17]),
        .Q(p_20_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[18]),
        .Q(p_21_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[19]),
        .Q(p_22_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[1]),
        .Q(p_2_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[20]),
        .Q(p_23_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[21]),
        .Q(p_24_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[22]),
        .Q(p_25_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[23]),
        .Q(p_26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[24]),
        .Q(p_27_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[25]),
        .Q(p_28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[26]),
        .Q(p_1_in26_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[27]),
        .Q(p_0_in28_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[28]),
        .Q(p_29_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[29]),
        .Q(p_30_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[2]),
        .Q(p_4_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[30]),
        .Q(p_31_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[31]),
        .Q(p_32_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[32]),
        .Q(p_33_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[33]),
        .Q(p_34_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[34]),
        .Q(p_35_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[35]),
        .Q(p_36_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[36]),
        .Q(p_3_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[3]),
        .Q(p_6_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[4]),
        .Q(p_7_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[5]),
        .Q(p_8_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[6]),
        .Q(p_9_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[7]),
        .Q(p_10_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[8]),
        .Q(p_11_in));
  FDCE #(
    .INIT(1'b0)) 
    \CASR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(p_0_in__0[9]),
        .Q(p_12_in));
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[0]_i_1 
       (.I0(seed_i[0]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[41] ),
        .O(\LFSR_reg[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[10]_i_1 
       (.I0(seed_i[10]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[9] ),
        .O(\LFSR_reg[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[11]_i_1 
       (.I0(seed_i[11]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[10] ),
        .O(\LFSR_reg[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[12]_i_1 
       (.I0(seed_i[12]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[11] ),
        .O(\LFSR_reg[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[13]_i_1 
       (.I0(seed_i[13]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[12] ),
        .O(\LFSR_reg[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[14]_i_1 
       (.I0(seed_i[14]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[13] ),
        .O(\LFSR_reg[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[15]_i_1 
       (.I0(seed_i[15]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[14] ),
        .O(\LFSR_reg[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[16]_i_1 
       (.I0(seed_i[16]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[15] ),
        .O(\LFSR_reg[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[17]_i_1 
       (.I0(seed_i[17]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[16] ),
        .O(\LFSR_reg[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[18]_i_1 
       (.I0(seed_i[18]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[17] ),
        .O(\LFSR_reg[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[19]_i_1 
       (.I0(seed_i[19]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[18] ),
        .O(\LFSR_reg[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[1]_i_1 
       (.I0(seed_i[1]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(\LFSR_reg_reg_n_0_[0] ),
        .O(\LFSR_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT4 #(
    .INIT(16'h8BB8)) 
    \LFSR_reg[20]_i_1 
       (.I0(seed_i[20]),
        .I1(loadseed_i),
        .I2(p_0_in),
        .I3(p_1_in0_in),
        .O(\LFSR_reg[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[21]_i_1 
       (.I0(seed_i[21]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[20] ),
        .O(\LFSR_reg[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[22]_i_1 
       (.I0(seed_i[22]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[21] ),
        .O(\LFSR_reg[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[23]_i_1 
       (.I0(seed_i[23]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[22] ),
        .O(\LFSR_reg[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[24]_i_1 
       (.I0(seed_i[24]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[23] ),
        .O(\LFSR_reg[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[25]_i_1 
       (.I0(seed_i[25]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[24] ),
        .O(\LFSR_reg[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[26]_i_1 
       (.I0(seed_i[26]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[25] ),
        .O(\LFSR_reg[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[27]_i_1 
       (.I0(seed_i[27]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[26] ),
        .O(\LFSR_reg[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[28]_i_1 
       (.I0(seed_i[28]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[27] ),
        .O(\LFSR_reg[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[29]_i_1 
       (.I0(seed_i[29]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[28] ),
        .O(\LFSR_reg[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[2]_i_1 
       (.I0(seed_i[2]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[1] ),
        .O(\LFSR_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[30]_i_1 
       (.I0(seed_i[30]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[29] ),
        .O(\LFSR_reg[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[31]_i_1 
       (.I0(seed_i[31]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[30] ),
        .O(\LFSR_reg[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[32]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[31] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[33]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[32] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[34]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[33] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[35]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[34] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[36]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[35] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[37]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[36] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[38]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[37] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[39]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[38] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[3]_i_1 
       (.I0(seed_i[3]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[2] ),
        .O(\LFSR_reg[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[40]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[39] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \LFSR_reg[41]_i_1 
       (.I0(p_1_in),
        .I1(p_0_in),
        .I2(loadseed_i),
        .O(\LFSR_reg[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \LFSR_reg[42]_i_1 
       (.I0(\LFSR_reg_reg_n_0_[41] ),
        .I1(loadseed_i),
        .O(\LFSR_reg[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[4]_i_1 
       (.I0(seed_i[4]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[3] ),
        .O(\LFSR_reg[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[5]_i_1 
       (.I0(seed_i[5]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[4] ),
        .O(\LFSR_reg[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[6]_i_1 
       (.I0(seed_i[6]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[5] ),
        .O(\LFSR_reg[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[7]_i_1 
       (.I0(seed_i[7]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[6] ),
        .O(\LFSR_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[8]_i_1 
       (.I0(seed_i[8]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[7] ),
        .O(\LFSR_reg[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \LFSR_reg[9]_i_1 
       (.I0(seed_i[9]),
        .I1(loadseed_i),
        .I2(\LFSR_reg_reg_n_0_[8] ),
        .O(\LFSR_reg[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \LFSR_reg_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .D(\LFSR_reg[0]_i_1_n_0 ),
        .PRE(\number_o[31]_i_2_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[10]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[11]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[12]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[13]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[14]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[15]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[16]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[17]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[18]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[19]_i_1_n_0 ),
        .Q(p_1_in0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[1]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[20]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[21]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[22]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[23]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[24]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[25]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[26]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[27]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[28]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[29]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[2]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[30]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[31]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[32] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[32]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[33] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[33]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[34] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[34]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[35] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[35]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[36] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[36]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[37] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[37]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[38] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[38]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[39] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[39]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[3]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[40] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[40]_i_1_n_0 ),
        .Q(p_1_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[41] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[41]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[42] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[42]_i_1_n_0 ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[4]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[5]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[6]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[7]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[8]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \LFSR_reg_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\LFSR_reg[9]_i_1_n_0 ),
        .Q(\LFSR_reg_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[0]_i_1 
       (.I0(\CASR_reg_reg_n_0_[0] ),
        .I1(\LFSR_reg_reg_n_0_[0] ),
        .O(\number_o[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[10]_i_1 
       (.I0(p_13_in),
        .I1(\LFSR_reg_reg_n_0_[10] ),
        .O(\number_o[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[11]_i_1 
       (.I0(p_14_in),
        .I1(\LFSR_reg_reg_n_0_[11] ),
        .O(\number_o[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[12]_i_1 
       (.I0(p_15_in),
        .I1(\LFSR_reg_reg_n_0_[12] ),
        .O(\number_o[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[13]_i_1 
       (.I0(p_16_in),
        .I1(\LFSR_reg_reg_n_0_[13] ),
        .O(\number_o[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[14]_i_1 
       (.I0(p_17_in),
        .I1(\LFSR_reg_reg_n_0_[14] ),
        .O(\number_o[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[15]_i_1 
       (.I0(p_18_in),
        .I1(\LFSR_reg_reg_n_0_[15] ),
        .O(\number_o[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[16]_i_1 
       (.I0(p_19_in),
        .I1(\LFSR_reg_reg_n_0_[16] ),
        .O(\number_o[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[17]_i_1 
       (.I0(p_20_in),
        .I1(\LFSR_reg_reg_n_0_[17] ),
        .O(\number_o[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[18]_i_1 
       (.I0(p_21_in),
        .I1(\LFSR_reg_reg_n_0_[18] ),
        .O(\number_o[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[19]_i_1 
       (.I0(p_22_in),
        .I1(p_1_in0_in),
        .O(\number_o[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[1]_i_1 
       (.I0(p_2_in),
        .I1(\LFSR_reg_reg_n_0_[1] ),
        .O(\number_o[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[20]_i_1 
       (.I0(p_23_in),
        .I1(\LFSR_reg_reg_n_0_[20] ),
        .O(\number_o[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[21]_i_1 
       (.I0(p_24_in),
        .I1(\LFSR_reg_reg_n_0_[21] ),
        .O(\number_o[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[22]_i_1 
       (.I0(p_25_in),
        .I1(\LFSR_reg_reg_n_0_[22] ),
        .O(\number_o[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[23]_i_1 
       (.I0(p_26_in),
        .I1(\LFSR_reg_reg_n_0_[23] ),
        .O(\number_o[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[24]_i_1 
       (.I0(p_27_in),
        .I1(\LFSR_reg_reg_n_0_[24] ),
        .O(\number_o[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[25]_i_1 
       (.I0(p_28_in),
        .I1(\LFSR_reg_reg_n_0_[25] ),
        .O(\number_o[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[26]_i_1 
       (.I0(p_1_in26_in),
        .I1(\LFSR_reg_reg_n_0_[26] ),
        .O(\number_o[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[27]_i_1 
       (.I0(p_0_in28_in),
        .I1(\LFSR_reg_reg_n_0_[27] ),
        .O(\number_o[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[28]_i_1 
       (.I0(p_29_in),
        .I1(\LFSR_reg_reg_n_0_[28] ),
        .O(\number_o[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[29]_i_1 
       (.I0(p_30_in),
        .I1(\LFSR_reg_reg_n_0_[29] ),
        .O(\number_o[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[2]_i_1 
       (.I0(p_4_in),
        .I1(\LFSR_reg_reg_n_0_[2] ),
        .O(\number_o[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[30]_i_1 
       (.I0(p_31_in),
        .I1(\LFSR_reg_reg_n_0_[30] ),
        .O(\number_o[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[31]_i_1 
       (.I0(p_32_in),
        .I1(\LFSR_reg_reg_n_0_[31] ),
        .O(\number_o[31]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \number_o[31]_i_2 
       (.I0(reset),
        .O(\number_o[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[3]_i_1 
       (.I0(p_6_in),
        .I1(\LFSR_reg_reg_n_0_[3] ),
        .O(\number_o[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[4]_i_1 
       (.I0(p_7_in),
        .I1(\LFSR_reg_reg_n_0_[4] ),
        .O(\number_o[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[5]_i_1 
       (.I0(p_8_in),
        .I1(\LFSR_reg_reg_n_0_[5] ),
        .O(\number_o[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[6]_i_1 
       (.I0(p_9_in),
        .I1(\LFSR_reg_reg_n_0_[6] ),
        .O(\number_o[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[7]_i_1 
       (.I0(p_10_in),
        .I1(\LFSR_reg_reg_n_0_[7] ),
        .O(\number_o[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[8]_i_1 
       (.I0(p_11_in),
        .I1(\LFSR_reg_reg_n_0_[8] ),
        .O(\number_o[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \number_o[9]_i_1 
       (.I0(p_12_in),
        .I1(\LFSR_reg_reg_n_0_[9] ),
        .O(\number_o[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[0] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[0]_i_1_n_0 ),
        .Q(number_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[10] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[10]_i_1_n_0 ),
        .Q(number_o[10]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[11] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[11]_i_1_n_0 ),
        .Q(number_o[11]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[12] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[12]_i_1_n_0 ),
        .Q(number_o[12]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[13] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[13]_i_1_n_0 ),
        .Q(number_o[13]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[14] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[14]_i_1_n_0 ),
        .Q(number_o[14]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[15] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[15]_i_1_n_0 ),
        .Q(number_o[15]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[16] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[16]_i_1_n_0 ),
        .Q(number_o[16]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[17] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[17]_i_1_n_0 ),
        .Q(number_o[17]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[18] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[18]_i_1_n_0 ),
        .Q(number_o[18]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[19] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[19]_i_1_n_0 ),
        .Q(number_o[19]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[1] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[1]_i_1_n_0 ),
        .Q(number_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[20] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[20]_i_1_n_0 ),
        .Q(number_o[20]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[21] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[21]_i_1_n_0 ),
        .Q(number_o[21]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[22] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[22]_i_1_n_0 ),
        .Q(number_o[22]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[23] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[23]_i_1_n_0 ),
        .Q(number_o[23]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[24] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[24]_i_1_n_0 ),
        .Q(number_o[24]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[25] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[25]_i_1_n_0 ),
        .Q(number_o[25]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[26] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[26]_i_1_n_0 ),
        .Q(number_o[26]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[27] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[27]_i_1_n_0 ),
        .Q(number_o[27]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[28] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[28]_i_1_n_0 ),
        .Q(number_o[28]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[29] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[29]_i_1_n_0 ),
        .Q(number_o[29]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[2] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[2]_i_1_n_0 ),
        .Q(number_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[30] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[30]_i_1_n_0 ),
        .Q(number_o[30]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[31] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[31]_i_1_n_0 ),
        .Q(number_o[31]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[3] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[3]_i_1_n_0 ),
        .Q(number_o[3]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[4] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[4]_i_1_n_0 ),
        .Q(number_o[4]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[5] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[5]_i_1_n_0 ),
        .Q(number_o[5]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[6] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[6]_i_1_n_0 ),
        .Q(number_o[6]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[7] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[7]_i_1_n_0 ),
        .Q(number_o[7]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[8] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[8]_i_1_n_0 ),
        .Q(number_o[8]));
  FDCE #(
    .INIT(1'b0)) 
    \number_o_reg[9] 
       (.C(clk),
        .CE(1'b1),
        .CLR(\number_o[31]_i_2_n_0 ),
        .D(\number_o[9]_i_1_n_0 ),
        .Q(number_o[9]));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench__1
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench__2
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench__3
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench__4
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench__5
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule

(* ORIG_REF_NAME = "s13207_bench" *) (* keep = "true" *) 
module switch_elements_s13207_bench__6
   (blif_clk_net,
    blif_reset_net,
    g43,
    g49,
    g633,
    g634,
    g635,
    g645,
    g647,
    g648,
    g690,
    g694,
    g698,
    g702,
    g722,
    g723,
    g751,
    g752,
    g753,
    g754,
    g755,
    g756,
    g757,
    g781,
    g941,
    g962,
    g1000,
    g1008,
    g1016,
    g1080,
    g1234,
    g1553,
    g1554,
    g206,
    g291,
    g372,
    g453,
    g534,
    g594,
    g785,
    g1006,
    g1015,
    g1017,
    g1246,
    g1724,
    g1783,
    g1798,
    g1804,
    g1810,
    g1817,
    g1824,
    g1829,
    g1870,
    g1871,
    g1894,
    g1911,
    g1944,
    g2662,
    g2844,
    g2888,
    g3077,
    g3096,
    g3130,
    g3159,
    g3191,
    g3829,
    g3859,
    g3860,
    g4267,
    g4316,
    g4370,
    g4371,
    g4372,
    g4373,
    g4655,
    g4657,
    g4660,
    g4661,
    g4663,
    g4664,
    g5143,
    g5164,
    g5571,
    g5669,
    g5678,
    g5682,
    g5684,
    g5687,
    g5729,
    g6207,
    g6212,
    g6223,
    g6236,
    g6269,
    g6425,
    g6648,
    g6653,
    g6675,
    g6849,
    g6850,
    g6895,
    g6909,
    g7048,
    g7063,
    g7103,
    g7283,
    g7284,
    g7285,
    g7286,
    g7287,
    g7288,
    g7289,
    g7290,
    g7291,
    g7292,
    g7293,
    g7294,
    g7295,
    g7298,
    g7423,
    g7424,
    g7425,
    g7474,
    g7504,
    g7505,
    g7506,
    g7507,
    g7508,
    g7514,
    g7729,
    g7730,
    g7731,
    g7732,
    g8216,
    g8217,
    g8218,
    g8219,
    g8234,
    g8661,
    g8663,
    g8872,
    g8958,
    g9128,
    g9132,
    g9204,
    g9280,
    g9297,
    g9299,
    g9305,
    g9308,
    g9310,
    g9312,
    g9314,
    g9378);
  input blif_clk_net;
  input blif_reset_net;
  input g43;
  input g49;
  input g633;
  input g634;
  input g635;
  input g645;
  input g647;
  input g648;
  input g690;
  input g694;
  input g698;
  input g702;
  input g722;
  input g723;
  input g751;
  input g752;
  input g753;
  input g754;
  input g755;
  input g756;
  input g757;
  input g781;
  input g941;
  input g962;
  input g1000;
  input g1008;
  input g1016;
  input g1080;
  input g1234;
  input g1553;
  input g1554;
  output g206;
  output g291;
  output g372;
  output g453;
  output g534;
  output g594;
  output g785;
  output g1006;
  output g1015;
  output g1017;
  output g1246;
  output g1724;
  output g1783;
  output g1798;
  output g1804;
  output g1810;
  output g1817;
  output g1824;
  output g1829;
  output g1870;
  output g1871;
  output g1894;
  output g1911;
  output g1944;
  output g2662;
  output g2844;
  output g2888;
  output g3077;
  output g3096;
  output g3130;
  output g3159;
  output g3191;
  output g3829;
  output g3859;
  output g3860;
  output g4267;
  output g4316;
  output g4370;
  output g4371;
  output g4372;
  output g4373;
  output g4655;
  output g4657;
  output g4660;
  output g4661;
  output g4663;
  output g4664;
  output g5143;
  output g5164;
  output g5571;
  output g5669;
  output g5678;
  output g5682;
  output g5684;
  output g5687;
  output g5729;
  output g6207;
  output g6212;
  output g6223;
  output g6236;
  output g6269;
  output g6425;
  output g6648;
  output g6653;
  output g6675;
  output g6849;
  output g6850;
  output g6895;
  output g6909;
  output g7048;
  output g7063;
  output g7103;
  output g7283;
  output g7284;
  output g7285;
  output g7286;
  output g7287;
  output g7288;
  output g7289;
  output g7290;
  output g7291;
  output g7292;
  output g7293;
  output g7294;
  output g7295;
  output g7298;
  output g7423;
  output g7424;
  output g7425;
  output g7474;
  output g7504;
  output g7505;
  output g7506;
  output g7507;
  output g7508;
  output g7514;
  output g7729;
  output g7730;
  output g7731;
  output g7732;
  output g8216;
  output g8217;
  output g8218;
  output g8219;
  output g8234;
  output g8661;
  output g8663;
  output g8872;
  output g8958;
  output g9128;
  output g9132;
  output g9204;
  output g9280;
  output g9297;
  output g9299;
  output g9305;
  output g9308;
  output g9310;
  output g9312;
  output g9314;
  output g9378;

  wire \<const0> ;
  wire blif_clk_net;
  wire blif_reset_net;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g10;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g100;
  wire g1000;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1004;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1005;
  wire g1006;
  wire g1006_INST_0_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1007;
  wire g1008;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1012;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1013;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1014;
  wire g1015;
  wire g1016;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1018;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1021;
  wire g1021_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1025;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1029;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g103;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1030;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1033;
  wire g1033_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1034;
  wire g1034_i_2_n_0;
  wire g1034_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1037;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g104;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1041;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1045;
  wire g1045_i_2_n_0;
  wire g1045_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1049;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g105;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1053;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1057;
  wire g1057_i_2_n_0;
  wire g1057_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1061;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1065;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1069;
  wire g1069_i_2_n_0;
  wire g1069_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1073;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1077;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g108;
  wire g1080;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1081;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1084;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1087;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g109;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1092;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1097;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g11;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g110;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1102;
  wire g1102_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1106;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1110;
  wire g1110_i_1_n_0;
  wire g1110_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1122;
  wire g1122_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1126;
  wire g1126_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g113;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1138;
  wire g1138_i_2_n_0;
  wire g1138_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g114;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1142;
  wire g1142_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1147;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1148;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1149;
  wire g1149_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1153;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1155;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1156;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1157;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1159;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1160;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1163;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1166;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1167;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g117;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1170;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1173;
  wire g1173_i_2_n_0;
  wire g1173_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1176;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g118;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1189;
  wire g1189_i_2_n_0;
  wire g1189_i_3_n_0;
  wire g1189_i_4_n_0;
  wire g1189_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1191;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1192;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1193;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1194;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1197;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1198;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g12;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1203;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1207;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g121;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1217;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g122;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1220;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1223;
  wire g1223_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1224;
  wire g1224_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1225;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1226;
  wire g1226_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1227;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1229;
  wire g1229_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1230;
  wire g1230_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1231;
  wire g1234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1244;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1245;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1247;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g125;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1250;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1251;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1253;
  wire g1253_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1254;
  wire g1254_i_2_n_0;
  wire g1254_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1257;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g126;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1260;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1263;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1266;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1267;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1268;
  wire g1268_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1269;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1271;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1272;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1276;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1280;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1284;
  wire g1284_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1288;
  wire g1288_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g129;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1296;
  wire g1296_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g13;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g130;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1300;
  wire g1300_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1304;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1307;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1308;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1310;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1311;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1319;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1320;
  wire g1320_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1322;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1323;
  wire g1323_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1324;
  wire g1324_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1325;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1326;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1327;
  wire g1327_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1328;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1329;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g133;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1330;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1333;
  wire g1333_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1339;
  wire g1339_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g134;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1345;
  wire g1345_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1348;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1351;
  wire g1351_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1354;
  wire g1354_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1357;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1360;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1363;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1364;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1366;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1369;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g137;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1370;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1372;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1379;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g138;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1380;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1381;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1382;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1383;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1384;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1385;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1386;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1388;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1389;
  wire g1389_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1391;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1392;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1399;
  wire g13_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1400;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1401;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1402;
  wire g1402_i_2_n_0;
  wire g1402_i_3_n_0;
  wire g1402_i_4_n_0;
  wire g1402_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1403;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1404;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1409;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g141;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1412;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1415;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1416;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g142;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1421;
  wire g1421_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1424;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1428;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1429;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1430;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1431;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1435;
  wire g1435_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1439;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1444;
  wire g1444_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1450;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1459;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g146;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1460;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1461;
  wire g1461_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1462;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1467;
  wire g1467_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1472;
  wire g1472_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1481;
  wire g1481_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1486;
  wire g1486_i_2_n_0;
  wire g1486_i_3_n_0;
  wire g1486_i_4_n_0;
  wire g1486_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1489;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1494;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1499;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g150;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1504;
  wire g1504_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1509;
  wire g1509_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1514;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1519;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g1524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1528;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1532;
  wire g1532_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1537;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g154;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1541;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1545;
  wire g1545_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g1549;
  wire g1549_i_2_n_0;
  wire g1553;
  wire g1554;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g158;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g16;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g162;
  wire g162_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g168;
  wire g1681;
  wire g1683;
  wire g1707;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g172;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g173;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g174;
  wire g1789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g179;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g180;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g181;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g182;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g183;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g184;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g185;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g186;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g190;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g195;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g196;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g199;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g2;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g20;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g200;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g201;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g202;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g205;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g207;
  wire g20_i_2_n_0;
  wire g20_i_3_n_0;
  wire g20_i_4_n_0;
  wire g20_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g21;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g210;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g211;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g212;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g213;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g214;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g215;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g216;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g219;
  wire g219_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g22;
  wire g2206;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g222;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g225;
  wire g2262;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g228;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g23;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g231;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g232;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g233;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g234;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g235;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g236;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g237;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g24;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g240;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g243;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g246;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g249;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g25;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g252;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g255;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g258;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g26;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g261;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g264;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g267;
  wire g267_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g27;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g270;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g273;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g274;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g275;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g278;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g28;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g281;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g284;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g29;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g290;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g292;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g293;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g294;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g295;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g296;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g297;
  wire g2_i_2_n_0;
  wire g2_i_3_n_0;
  wire g2_i_4_n_0;
  wire g2_i_5_n_0;
  wire g2_i_6_n_0;
  wire g2_i_7_n_0;
  (* RTL_KEEP = "true" *) wire g3;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g30;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g300;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g303;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g306;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g31;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g312;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g313;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g314;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g315;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g316;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g317;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g318;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g32;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g321;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g324;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g327;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g33;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g330;
  wire g330_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g333;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g336;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g339;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g342;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g345;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g348;
  wire g348_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g351;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g354;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g355;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g356;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g359;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g362;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g365;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g368;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g37;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g371;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g373;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g374;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g375;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g376;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g377;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g378;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g38;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g381;
  wire g381_i_1_n_0;
  wire g3832;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g384;
  wire g3863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g387;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g390;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g393;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g394;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g395;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g396;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g397;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g398;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g399;
  (* RTL_KEEP = "true" *) wire g4;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g402;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g405;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g408;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g41;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g411;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g414;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g417;
  (* RTL_KEEP = "true" *) wire g42;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g420;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g423;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g426;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g429;
  wire g43;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g432;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g435;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g436;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g437;
  (* RTL_KEEP = "true" *) wire g44;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g440;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g443;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g446;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g449;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g45;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g452;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g454;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g455;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g456;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g457;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g458;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g459;
  wire g4598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g46;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g462;
  wire g462_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g465;
  wire g4652;
  wire g4654;
  wire g4655;
  wire g4656;
  wire g4657;
  wire g4657_INST_0_i_1_n_0;
  wire g4658;
  wire g4660;
  wire g4661;
  wire g4663;
  wire g4664;
  wire g4665;
  wire g4666;
  wire g4668;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g468;
  wire g4681;
  (* RTL_KEEP = "true" *) wire g47;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g471;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g474;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g475;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g476;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g477;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g478;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g479;
  wire g4792;
  wire g47_i_2_n_0;
  wire g47_i_3_n_0;
  wire g47_i_4_n_0;
  wire g47_i_5_n_0;
  wire g47_i_6_n_0;
  wire g47_i_7_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g48;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g480;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g483;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g486;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g489;
  wire g49;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g492;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g495;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g498;
  wire g498_i_1_n_0;
  wire g498_i_2_n_0;
  wire g4_i_2_n_0;
  wire g4_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g5;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g501;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g504;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g507;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g510;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g513;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g516;
  wire g5163;
  wire g5164;
  wire g5165;
  wire g5166;
  wire g5167;
  wire g5168;
  wire g5169;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g517;
  wire g5170;
  wire g5172;
  wire g5173;
  wire g5174;
  wire g5175;
  wire g5177;
  wire g5178;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g518;
  wire g5180;
  wire g5182;
  wire g5183;
  wire g5184;
  wire g5186;
  wire g5187;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g52;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g521;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g524;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g527;
  wire g5287;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g530;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g533;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g535;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g536;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g539;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g540;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g543;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g544;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g547;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g55;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g550;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g553;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g556;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g557;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g560;
  wire g560_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g563;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g566;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g567;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g570;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g573;
  wire g5730;
  wire g5731;
  wire g5732;
  wire g5733;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5737;
  wire g5738;
  wire g5739;
  wire g573_i_1_n_0;
  wire g573_i_2_n_0;
  wire g5740;
  wire g5742;
  wire g5743;
  wire g5744;
  wire g5745;
  wire g5746;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g576;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g579;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g58;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g580;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g583;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g584;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g587;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g588;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g591;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g595;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g596;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g597;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g598;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g599;
  (* RTL_KEEP = "true" *) wire g6;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g600;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g601;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g602;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g603;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g604;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g605;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g606;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g607;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g608;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g609;
  wire g6098;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g610;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g611;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g612;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g613;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g614;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g615;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g616;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g617;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g618;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g619;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g62;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g620;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g621;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g622;
  wire g6223;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g623;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g624;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g625;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g626;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g627;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g628;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g629;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g630;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g631;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g632;
  wire g633;
  wire g634;
  wire g635;
  wire g6371;
  wire g6372;
  wire g6377;
  wire g6378;
  wire g6379;
  wire g6380;
  wire g6381;
  wire g6382;
  wire g6383;
  wire g6384;
  wire g6385;
  wire g6386;
  wire g6391;
  wire g6392;
  wire g645;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g646;
  wire g647;
  wire g648;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g65;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g652;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g661;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g665;
  wire g6664;
  wire g6675;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g669;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g673;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g677;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g68;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g681;
  wire g6849;
  wire g6849_INST_0_i_1_n_0;
  wire g6849_INST_0_i_2_n_0;
  wire g6849_INST_0_i_3_n_0;
  wire g6849_INST_0_i_4_n_0;
  wire g6849_INST_0_i_5_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g685;
  wire g6850;
  wire g6852;
  wire g6853;
  wire g6854;
  wire g6856;
  wire g6857;
  wire g6858;
  wire g6859;
  wire g6861;
  wire g6862;
  wire g6864;
  wire g6866;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6870;
  wire g6871;
  wire g6872;
  wire g6873;
  wire g6874;
  wire g6875;
  wire g6876;
  wire g6877;
  wire g6878;
  wire g6879;
  wire g6880;
  wire g6881;
  wire g6882;
  wire g6883;
  wire g6884;
  wire g6885;
  wire g6886;
  wire g6887;
  wire g6888;
  wire g6889;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g689;
  wire g6890;
  wire g6891;
  wire g6895;
  wire g689_i_2_n_0;
  wire g689_i_3_n_0;
  wire g689_i_4_n_0;
  wire g689_i_5_n_0;
  wire g689_i_6_n_0;
  wire g690;
  wire g694;
  wire g698;
  (* RTL_KEEP = "true" *) wire g7;
  wire g702;
  wire g7048;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g706;
  wire g706_i_1_n_0;
  wire g706_i_2_n_0;
  wire g7099;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g71;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g710;
  wire g7100;
  wire g7101;
  wire g7102;
  wire g7103;
  wire g7103_INST_0_i_1_n_0;
  wire g7103_INST_0_i_2_n_0;
  wire g7105;
  wire g7106;
  wire g7107;
  wire g7108;
  wire g7109;
  wire g7110;
  wire g7111;
  wire g7112;
  wire g7113;
  wire g7114;
  wire g7115;
  wire g7116;
  wire g7117;
  wire g7118;
  wire g7119;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g714;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g718;
  wire g7217;
  wire g722;
  wire g723;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g727;
  wire g7283;
  wire g7283_INST_0_i_1_n_0;
  wire g7283_INST_0_i_2_n_0;
  wire g7284;
  wire g7285;
  wire g7286;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7291_INST_0_i_1_n_0;
  wire g7292;
  wire g7293;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g730;
  wire g7300;
  wire g7302;
  wire g7303;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g734;
  wire g734_i_1_n_0;
  wire g7367;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g74;
  wire g7406;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g741;
  wire g741_i_2_n_0;
  wire g741_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g746;
  wire g746_i_2_n_0;
  wire g7474;
  wire g7480;
  wire g751;
  wire g7510;
  wire g7511;
  wire g7514;
  wire g7515;
  wire g7516;
  wire g7518;
  wire g7519;
  wire g752;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7523;
  wire g7524;
  wire g7525;
  wire g7527;
  wire g7528;
  wire g7529;
  wire g753;
  wire g754;
  wire g755;
  wire g756;
  wire g7566;
  wire g757;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g758;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g759;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g760;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g761;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g762;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g763;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g764;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g765;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g766;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g767;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g768;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g769;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g77;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g770;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g771;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g772;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g773;
  wire g7731;
  wire g7739;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g774;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g775;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g775_i_2_n_0;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g778;
  wire g7780;
  wire g7781;
  wire g778_i_2_n_0;
  wire g781;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g782;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g786;
  wire g786_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g789;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g792;
  wire g792_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g795;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g799;
  wire g799_i_2_n_0;
  (* RTL_KEEP = "true" *) wire g8;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g80;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g803;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g806;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g809;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g812;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g815;
  wire g815_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g819;
  wire g819_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g822;
  wire g8220;
  wire g8221;
  wire g8222;
  wire g8224;
  wire g8226;
  wire g8227;
  wire g8228;
  wire g822_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g825;
  wire g825_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g828;
  wire g828_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g83;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g831;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g834;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g837;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g840;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g843;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g846;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g849;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g852;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g855;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g859;
  wire g859_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g86;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g863;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g866;
  wire g8663;
  wire g8664;
  wire g8665;
  wire g8666;
  wire g8667;
  wire g8668;
  wire g8669;
  wire g8670;
  wire g8671;
  wire g8673;
  wire g8674;
  wire g8675;
  wire g8676;
  wire g8677;
  wire g8678;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g871;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g874;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g875;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g878;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g883;
  wire g8865;
  wire g8867;
  wire g8869;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g887;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8872_INST_0_i_1_n_0;
  wire g8873;
  wire g8875;
  wire g887_i_2_n_0;
  wire g887_i_3_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g888;
  wire g888_i_2_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g889;
  wire g889_i_2_n_0;
  wire g889_i_3_n_0;
  wire g889_i_4_n_0;
  wire g889_i_5_n_0;
  wire g889_i_6_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g89;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g890;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g891;
  wire g8956;
  wire g8957;
  wire g8958;
  wire g8959;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g896;
  wire g8960;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g9;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g901;
  wire g9034;
  wire g9035;
  wire g9036;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g906;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g911;
  wire g9117;
  wire g9132;
  wire g9133;
  wire g9134;
  wire g9145;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g916;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g92;
  wire g9204;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g921;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g926;
  wire g9280;
  wire g9280_INST_0_i_10_n_0;
  wire g9280_INST_0_i_11_n_0;
  wire g9280_INST_0_i_12_n_0;
  wire g9280_INST_0_i_13_n_0;
  wire g9280_INST_0_i_14_n_0;
  wire g9280_INST_0_i_15_n_0;
  wire g9280_INST_0_i_16_n_0;
  wire g9280_INST_0_i_17_n_0;
  wire g9280_INST_0_i_18_n_0;
  wire g9280_INST_0_i_19_n_0;
  wire g9280_INST_0_i_1_n_0;
  wire g9280_INST_0_i_20_n_0;
  wire g9280_INST_0_i_21_n_0;
  wire g9280_INST_0_i_22_n_0;
  wire g9280_INST_0_i_23_n_0;
  wire g9280_INST_0_i_24_n_0;
  wire g9280_INST_0_i_25_n_0;
  wire g9280_INST_0_i_26_n_0;
  wire g9280_INST_0_i_27_n_0;
  wire g9280_INST_0_i_28_n_0;
  wire g9280_INST_0_i_29_n_0;
  wire g9280_INST_0_i_2_n_0;
  wire g9280_INST_0_i_30_n_0;
  wire g9280_INST_0_i_31_n_0;
  wire g9280_INST_0_i_32_n_0;
  wire g9280_INST_0_i_33_n_0;
  wire g9280_INST_0_i_34_n_0;
  wire g9280_INST_0_i_35_n_0;
  wire g9280_INST_0_i_36_n_0;
  wire g9280_INST_0_i_3_n_0;
  wire g9280_INST_0_i_4_n_0;
  wire g9280_INST_0_i_5_n_0;
  wire g9280_INST_0_i_6_n_0;
  wire g9280_INST_0_i_7_n_0;
  wire g9280_INST_0_i_8_n_0;
  wire g9280_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g929;
  wire g9297;
  wire g9297_INST_0_i_10_n_0;
  wire g9297_INST_0_i_11_n_0;
  wire g9297_INST_0_i_12_n_0;
  wire g9297_INST_0_i_13_n_0;
  wire g9297_INST_0_i_14_n_0;
  wire g9297_INST_0_i_15_n_0;
  wire g9297_INST_0_i_16_n_0;
  wire g9297_INST_0_i_17_n_0;
  wire g9297_INST_0_i_18_n_0;
  wire g9297_INST_0_i_19_n_0;
  wire g9297_INST_0_i_20_n_0;
  wire g9297_INST_0_i_21_n_0;
  wire g9297_INST_0_i_22_n_0;
  wire g9297_INST_0_i_23_n_0;
  wire g9297_INST_0_i_24_n_0;
  wire g9297_INST_0_i_2_n_0;
  wire g9297_INST_0_i_3_n_0;
  wire g9297_INST_0_i_4_n_0;
  wire g9297_INST_0_i_5_n_0;
  wire g9297_INST_0_i_6_n_0;
  wire g9297_INST_0_i_7_n_0;
  wire g9297_INST_0_i_8_n_0;
  wire g9297_INST_0_i_9_n_0;
  wire g9299;
  wire g9299_INST_0_i_10_n_0;
  wire g9299_INST_0_i_11_n_0;
  wire g9299_INST_0_i_12_n_0;
  wire g9299_INST_0_i_13_n_0;
  wire g9299_INST_0_i_14_n_0;
  wire g9299_INST_0_i_15_n_0;
  wire g9299_INST_0_i_16_n_0;
  wire g9299_INST_0_i_17_n_0;
  wire g9299_INST_0_i_18_n_0;
  wire g9299_INST_0_i_19_n_0;
  wire g9299_INST_0_i_1_n_0;
  wire g9299_INST_0_i_20_n_0;
  wire g9299_INST_0_i_21_n_0;
  wire g9299_INST_0_i_22_n_0;
  wire g9299_INST_0_i_23_n_0;
  wire g9299_INST_0_i_24_n_0;
  wire g9299_INST_0_i_25_n_0;
  wire g9299_INST_0_i_26_n_0;
  wire g9299_INST_0_i_27_n_0;
  wire g9299_INST_0_i_28_n_0;
  wire g9299_INST_0_i_29_n_0;
  wire g9299_INST_0_i_2_n_0;
  wire g9299_INST_0_i_30_n_0;
  wire g9299_INST_0_i_31_n_0;
  wire g9299_INST_0_i_32_n_0;
  wire g9299_INST_0_i_3_n_0;
  wire g9299_INST_0_i_4_n_0;
  wire g9299_INST_0_i_5_n_0;
  wire g9299_INST_0_i_6_n_0;
  wire g9299_INST_0_i_7_n_0;
  wire g9299_INST_0_i_8_n_0;
  wire g9299_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g93;
  wire g9305;
  wire g9305_INST_0_i_10_n_0;
  wire g9305_INST_0_i_11_n_0;
  wire g9305_INST_0_i_12_n_0;
  wire g9305_INST_0_i_13_n_0;
  wire g9305_INST_0_i_14_n_0;
  wire g9305_INST_0_i_15_n_0;
  wire g9305_INST_0_i_16_n_0;
  wire g9305_INST_0_i_17_n_0;
  wire g9305_INST_0_i_18_n_0;
  wire g9305_INST_0_i_19_n_0;
  wire g9305_INST_0_i_1_n_0;
  wire g9305_INST_0_i_20_n_0;
  wire g9305_INST_0_i_21_n_0;
  wire g9305_INST_0_i_22_n_0;
  wire g9305_INST_0_i_23_n_0;
  wire g9305_INST_0_i_24_n_0;
  wire g9305_INST_0_i_25_n_0;
  wire g9305_INST_0_i_26_n_0;
  wire g9305_INST_0_i_27_n_0;
  wire g9305_INST_0_i_28_n_0;
  wire g9305_INST_0_i_29_n_0;
  wire g9305_INST_0_i_2_n_0;
  wire g9305_INST_0_i_30_n_0;
  wire g9305_INST_0_i_31_n_0;
  wire g9305_INST_0_i_32_n_0;
  wire g9305_INST_0_i_33_n_0;
  wire g9305_INST_0_i_3_n_0;
  wire g9305_INST_0_i_4_n_0;
  wire g9305_INST_0_i_5_n_0;
  wire g9305_INST_0_i_6_n_0;
  wire g9305_INST_0_i_7_n_0;
  wire g9305_INST_0_i_8_n_0;
  wire g9305_INST_0_i_9_n_0;
  wire g9308;
  wire g9308_INST_0_i_10_n_0;
  wire g9308_INST_0_i_11_n_0;
  wire g9308_INST_0_i_12_n_0;
  wire g9308_INST_0_i_13_n_0;
  wire g9308_INST_0_i_14_n_0;
  wire g9308_INST_0_i_15_n_0;
  wire g9308_INST_0_i_16_n_0;
  wire g9308_INST_0_i_17_n_0;
  wire g9308_INST_0_i_18_n_0;
  wire g9308_INST_0_i_19_n_0;
  wire g9308_INST_0_i_1_n_0;
  wire g9308_INST_0_i_20_n_0;
  wire g9308_INST_0_i_21_n_0;
  wire g9308_INST_0_i_22_n_0;
  wire g9308_INST_0_i_23_n_0;
  wire g9308_INST_0_i_24_n_0;
  wire g9308_INST_0_i_2_n_0;
  wire g9308_INST_0_i_3_n_0;
  wire g9308_INST_0_i_4_n_0;
  wire g9308_INST_0_i_5_n_0;
  wire g9308_INST_0_i_6_n_0;
  wire g9308_INST_0_i_7_n_0;
  wire g9308_INST_0_i_8_n_0;
  wire g9308_INST_0_i_9_n_0;
  wire g9310;
  wire g9310_INST_0_i_10_n_0;
  wire g9310_INST_0_i_11_n_0;
  wire g9310_INST_0_i_12_n_0;
  wire g9310_INST_0_i_13_n_0;
  wire g9310_INST_0_i_14_n_0;
  wire g9310_INST_0_i_1_n_0;
  wire g9310_INST_0_i_2_n_0;
  wire g9310_INST_0_i_3_n_0;
  wire g9310_INST_0_i_4_n_0;
  wire g9310_INST_0_i_5_n_0;
  wire g9310_INST_0_i_6_n_0;
  wire g9310_INST_0_i_7_n_0;
  wire g9310_INST_0_i_8_n_0;
  wire g9310_INST_0_i_9_n_0;
  wire g9312;
  wire g9312_INST_0_i_10_n_0;
  wire g9312_INST_0_i_11_n_0;
  wire g9312_INST_0_i_12_n_0;
  wire g9312_INST_0_i_1_n_0;
  wire g9312_INST_0_i_2_n_0;
  wire g9312_INST_0_i_3_n_0;
  wire g9312_INST_0_i_4_n_0;
  wire g9312_INST_0_i_5_n_0;
  wire g9312_INST_0_i_6_n_0;
  wire g9312_INST_0_i_7_n_0;
  wire g9312_INST_0_i_8_n_0;
  wire g9312_INST_0_i_9_n_0;
  wire g9314;
  wire g9314_INST_0_i_10_n_0;
  wire g9314_INST_0_i_11_n_0;
  wire g9314_INST_0_i_2_n_0;
  wire g9314_INST_0_i_3_n_0;
  wire g9314_INST_0_i_4_n_0;
  wire g9314_INST_0_i_5_n_0;
  wire g9314_INST_0_i_6_n_0;
  wire g9314_INST_0_i_7_n_0;
  wire g9314_INST_0_i_8_n_0;
  wire g9314_INST_0_i_9_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g933;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g936;
  wire g9360;
  wire g9361;
  wire g9362;
  wire g9372;
  wire g9373;
  wire g9374;
  wire g9375;
  wire g9376;
  wire g9378;
  wire g9378_INST_0_i_10_n_0;
  wire g9378_INST_0_i_11_n_0;
  wire g9378_INST_0_i_12_n_0;
  wire g9378_INST_0_i_13_n_0;
  wire g9378_INST_0_i_14_n_0;
  wire g9378_INST_0_i_15_n_0;
  wire g9378_INST_0_i_16_n_0;
  wire g9378_INST_0_i_17_n_0;
  wire g9378_INST_0_i_18_n_0;
  wire g9378_INST_0_i_19_n_0;
  wire g9378_INST_0_i_20_n_0;
  wire g9378_INST_0_i_21_n_0;
  wire g9378_INST_0_i_22_n_0;
  wire g9378_INST_0_i_23_n_0;
  wire g9378_INST_0_i_24_n_0;
  wire g9378_INST_0_i_25_n_0;
  wire g9378_INST_0_i_26_n_0;
  wire g9378_INST_0_i_27_n_0;
  wire g9378_INST_0_i_28_n_0;
  wire g9378_INST_0_i_29_n_0;
  wire g9378_INST_0_i_2_n_0;
  wire g9378_INST_0_i_30_n_0;
  wire g9378_INST_0_i_31_n_0;
  wire g9378_INST_0_i_32_n_0;
  wire g9378_INST_0_i_33_n_0;
  wire g9378_INST_0_i_3_n_0;
  wire g9378_INST_0_i_4_n_0;
  wire g9378_INST_0_i_5_n_0;
  wire g9378_INST_0_i_6_n_0;
  wire g9378_INST_0_i_7_n_0;
  wire g9378_INST_0_i_8_n_0;
  wire g9378_INST_0_i_9_n_0;
  wire g9386;
  wire g9389;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g94;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g940;
  wire g941;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g942;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g943;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g944;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g945;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g948;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g949;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g95;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g950;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g951;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g952;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g953;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g954;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g955;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g959;
  wire g962;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g963;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g966;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g969;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g970;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g971;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g972;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g973;
  wire g973_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g976;
  wire g976_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g979;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g98;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g984;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g985;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* S *) 
  (* shreg_extract = "no" *) wire g99;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g990;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g995;
  wire g995_i_1_n_0;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g998;
  (* DONT_TOUCH *) (* RTL_KEEP = "true" *) (* shreg_extract = "no" *) wire g999;

  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g206 = g1460;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g291 = g1460;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g372 = g1460;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g453 = g1460;
  assign g5143 = g1554;
  assign g534 = g1460;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g594 = g1460;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6236 = g7731;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7063 = g8663;
  assign g7294 = g7295;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7732 = g6223;
  assign g785 = g888;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = g6675;
  assign g8234 = g9132;
  assign g8661 = \<const0> ;
  assign g9128 = g9204;
  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h2)) 
    g1004_i_1
       (.I0(g43),
        .I1(g162),
        .O(g7105));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1004_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7105),
        .Q(g1004));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1005_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1004),
        .Q(g1005));
  LUT4 #(
    .INIT(16'h0800)) 
    g1006_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g162),
        .I2(g1000),
        .I3(g43),
        .O(g1006));
  LUT6 #(
    .INIT(64'h0000020002000200)) 
    g1006_INST_0_i_1
       (.I0(g8872_INST_0_i_1_n_0),
        .I1(g979),
        .I2(g1034),
        .I3(g7103_INST_0_i_1_n_0),
        .I4(g976),
        .I5(g43),
        .O(g1006_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g1007_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g43),
        .I3(g10),
        .I4(g1),
        .I5(g162),
        .O(g8867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1007_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8867),
        .Q(g1007));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g100_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g99),
        .Q(g100));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1012_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g43),
        .Q(g1012));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1013_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1014),
        .Q(g1013));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1014_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1012),
        .Q(g1014));
  LUT4 #(
    .INIT(16'h8000)) 
    g1015_INST_0
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1013),
        .I2(g162),
        .I3(g1),
        .O(g1015));
  LUT5 #(
    .INIT(32'h0000FF54)) 
    g1018_i_1
       (.I0(g1018),
        .I1(g1025),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1018_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8869),
        .Q(g1018));
  LUT5 #(
    .INIT(32'h00000098)) 
    g1021_i_1
       (.I0(g1018),
        .I1(g1021),
        .I2(g1025),
        .I3(g1021_i_2_n_0),
        .I4(g1029),
        .O(g8870));
  LUT4 #(
    .INIT(16'h0DFF)) 
    g1021_i_2
       (.I0(g1033),
        .I1(g1029),
        .I2(g1034),
        .I3(g43),
        .O(g1021_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1021_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8870),
        .Q(g1021));
  LUT5 #(
    .INIT(32'h0000FFA8)) 
    g1025_i_1
       (.I0(g1025),
        .I1(g1018),
        .I2(g1021),
        .I3(g1029),
        .I4(g1021_i_2_n_0),
        .O(g8871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1025_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8871),
        .Q(g1025));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1029_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g168),
        .Q(g1029));
  LUT5 #(
    .INIT(32'h00000800)) 
    g1030_i_1
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .I3(g1034),
        .I4(g146),
        .O(g7518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1030_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7518),
        .Q(g1030));
  LUT6 #(
    .INIT(64'h4444445455555555)) 
    g1033_i_1
       (.I0(g7406),
        .I1(g1033_i_2_n_0),
        .I2(g1018),
        .I3(g1021),
        .I4(g1025),
        .I5(g1034_i_2_n_0),
        .O(g9034));
  LUT3 #(
    .INIT(8'h40)) 
    g1033_i_2
       (.I0(g1029),
        .I1(g1033),
        .I2(g43),
        .O(g1033_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1033_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9034),
        .Q(g1033));
  LUT5 #(
    .INIT(32'hFD00FDFD)) 
    g1034_i_1
       (.I0(g995),
        .I1(g985),
        .I2(g990),
        .I3(g1034),
        .I4(g1034_i_2_n_0),
        .O(g8957));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    g1034_i_2
       (.I0(g7566),
        .I1(g1034_i_3_n_0),
        .I2(g999),
        .I3(g1000),
        .I4(g998),
        .I5(g1),
        .O(g1034_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    g1034_i_3
       (.I0(g1),
        .I1(g10),
        .I2(g43),
        .I3(g1008),
        .I4(g1007),
        .I5(g1016),
        .O(g1034_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1034_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8957),
        .Q(g1034));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1037_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149),
        .I3(g1149_i_2_n_0),
        .I4(g1037),
        .O(g7519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1037_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7519),
        .Q(g1037));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g103_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g100),
        .Q(g103));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1041_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .I4(g1037),
        .I5(g1041),
        .O(g7765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1041_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7765),
        .Q(g1041));
  LUT4 #(
    .INIT(16'h7007)) 
    g1045_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .O(g8224));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    g1045_i_2
       (.I0(g1037),
        .I1(g1149),
        .I2(g1041),
        .I3(g1045_i_3_n_0),
        .I4(g1251),
        .I5(g1158),
        .O(g1045_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1045_i_3
       (.I0(g1134),
        .I1(g1130),
        .I2(g1138),
        .I3(g1092),
        .O(g1045_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1045_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8224),
        .Q(g1045));
  LUT5 #(
    .INIT(32'h77070070)) 
    g1049_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045),
        .I3(g1045_i_2_n_0),
        .I4(g1049),
        .O(g8673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1049_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8673),
        .Q(g1049));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g104_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g104));
  LUT6 #(
    .INIT(64'h7077777707000000)) 
    g1053_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1045_i_2_n_0),
        .I3(g1045),
        .I4(g1049),
        .I5(g1053),
        .O(g8873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1053_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8873),
        .Q(g1053));
  LUT4 #(
    .INIT(16'h0770)) 
    g1057_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .O(g8959));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    g1057_i_2
       (.I0(g1251),
        .I1(g1158),
        .I2(g1049),
        .I3(g1045),
        .I4(g1053),
        .I5(g1057_i_3_n_0),
        .O(g1057_i_2_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g1057_i_3
       (.I0(g1045_i_3_n_0),
        .I1(g1041),
        .I2(g1149),
        .I3(g1037),
        .O(g1057_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1057_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8959),
        .Q(g1057));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g105_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g104),
        .Q(g105));
  LUT5 #(
    .INIT(32'h07777000)) 
    g1061_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1057_i_2_n_0),
        .I3(g1057),
        .I4(g1061),
        .O(g9035));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1061_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9035),
        .Q(g1061));
  LUT6 #(
    .INIT(64'h0777777770000000)) 
    g1065_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1061),
        .I3(g1057),
        .I4(g1057_i_2_n_0),
        .I5(g1065),
        .O(g9117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1065_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9117),
        .Q(g1065));
  LUT4 #(
    .INIT(16'h0770)) 
    g1069_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069),
        .I3(g1069_i_2_n_0),
        .O(g9134));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1069_i_2
       (.I0(g1065),
        .I1(g1061),
        .I2(g1069_i_3_n_0),
        .I3(g1049),
        .I4(g1053),
        .I5(g1057),
        .O(g1069_i_2_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1069_i_3
       (.I0(g1045),
        .I1(g1138_i_3_n_0),
        .I2(g1045_i_3_n_0),
        .I3(g1041),
        .I4(g1149),
        .I5(g1037),
        .O(g1069_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1069_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9134),
        .Q(g1069));
  LUT4 #(
    .INIT(16'h7444)) 
    g1073_i_1
       (.I0(g1158),
        .I1(g1073),
        .I2(g1069_i_2_n_0),
        .I3(g1069),
        .O(g9145));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1073_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9145),
        .Q(g1073));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1077_i_1
       (.I0(g7217),
        .I1(g1167),
        .I2(g1173),
        .I3(g1166),
        .I4(g1170),
        .O(g7767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1077_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7767),
        .Q(g1077));
  LUT3 #(
    .INIT(8'h3A)) 
    g1081_i_1
       (.I0(g1080),
        .I1(g1176),
        .I2(g1081),
        .O(g6852));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1081_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6852),
        .Q(g1081));
  LUT5 #(
    .INIT(32'h00807F80)) 
    g1084_i_1
       (.I0(g1179),
        .I1(g652),
        .I2(g1158),
        .I3(g1084),
        .I4(g1077),
        .O(g7106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1084_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7106),
        .Q(g1084));
  LUT3 #(
    .INIT(8'h06)) 
    g1087_i_1
       (.I0(g1148),
        .I1(g1087),
        .I2(g1097),
        .O(g6853));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1087_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6853),
        .Q(g1087));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g108_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g105),
        .Q(g108));
  LUT4 #(
    .INIT(16'h7304)) 
    g1092_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1251),
        .I3(g1092),
        .O(g7520));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1092_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7520),
        .Q(g1092));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1097_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1185),
        .Q(g1097));
  LUT4 #(
    .INIT(16'h006A)) 
    g1098_i_1
       (.I0(g1098),
        .I1(g1148),
        .I2(g1087),
        .I3(g1097),
        .O(g6854));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1098_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6854),
        .Q(g1098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g109_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g10_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g10));
  LUT5 #(
    .INIT(32'h15554000)) 
    g1102_i_1
       (.I0(g1097),
        .I1(g1087),
        .I2(g1098),
        .I3(g1148),
        .I4(g1102),
        .O(g1102_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1102_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1102_i_1_n_0),
        .Q(g1102));
  LUT6 #(
    .INIT(64'hBEEEEEEEEEEEEEEE)) 
    g1106_i_1
       (.I0(g1097),
        .I1(g1106),
        .I2(g1148),
        .I3(g1102),
        .I4(g1087),
        .I5(g1098),
        .O(g7107));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1106_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7107),
        .Q(g1106));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g109),
        .Q(g110));
  LUT3 #(
    .INIT(8'hEB)) 
    g1110_i_1
       (.I0(g1097),
        .I1(g1110_i_2_n_0),
        .I2(g1110),
        .O(g1110_i_1_n_0));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g1110_i_2
       (.I0(g1102),
        .I1(g1106),
        .I2(g1098),
        .I3(g1087),
        .I4(g1148),
        .O(g1110_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1110_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1110_i_1_n_0),
        .Q(g1110));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1114_i_1
       (.I0(g1097),
        .I1(g1110),
        .I2(g1110_i_2_n_0),
        .I3(g1114),
        .O(g7521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7521),
        .Q(g1114));
  LUT5 #(
    .INIT(32'hFFAABFEA)) 
    g1118_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .O(g7766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7766),
        .Q(g1118));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAEAAA)) 
    g1122_i_1
       (.I0(g1097),
        .I1(g1114),
        .I2(g1110),
        .I3(g1118),
        .I4(g1110_i_2_n_0),
        .I5(g1122),
        .O(g1122_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1122_i_1_n_0),
        .Q(g1122));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1126_i_1
       (.I0(g1097),
        .I1(g1122),
        .I2(g1126_i_2_n_0),
        .I3(g1126),
        .O(g8674));
  LUT4 #(
    .INIT(16'hFF7F)) 
    g1126_i_2
       (.I0(g1114),
        .I1(g1110),
        .I2(g1118),
        .I3(g1110_i_2_n_0),
        .O(g1126_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8674),
        .Q(g1126));
  LUT5 #(
    .INIT(32'h4F5F1000)) 
    g1130_i_1
       (.I0(g1073),
        .I1(g1251),
        .I2(g1158),
        .I3(g1092),
        .I4(g1130),
        .O(g7522));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7522),
        .Q(g1130));
  LUT6 #(
    .INIT(64'h55FF15FF00004000)) 
    g1134_i_1
       (.I0(g1073),
        .I1(g1130),
        .I2(g1092),
        .I3(g1158),
        .I4(g1251),
        .I5(g1134),
        .O(g7523));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7523),
        .Q(g1134));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1138_i_1
       (.I0(g1138_i_2_n_0),
        .I1(g1134),
        .I2(g1138_i_3_n_0),
        .I3(g1092),
        .I4(g1130),
        .I5(g1138),
        .O(g7524));
  LUT2 #(
    .INIT(4'h7)) 
    g1138_i_2
       (.I0(g1158),
        .I1(g1073),
        .O(g1138_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g1138_i_3
       (.I0(g1158),
        .I1(g1251),
        .O(g1138_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7524),
        .Q(g1138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g113_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g110),
        .Q(g113));
  LUT5 #(
    .INIT(32'h51550400)) 
    g1142_i_1
       (.I0(g1097),
        .I1(g1126),
        .I2(g1126_i_2_n_0),
        .I3(g1122),
        .I4(g1142),
        .O(g1142_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1142_i_1_n_0),
        .Q(g1142));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1146_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1084),
        .Q(g1146));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1147_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1146),
        .Q(g1147));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1148_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1147),
        .Q(g1148));
  LUT4 #(
    .INIT(16'h7007)) 
    g1149_i_1
       (.I0(g1073),
        .I1(g1158),
        .I2(g1149_i_2_n_0),
        .I3(g1149),
        .O(g7525));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1149_i_2
       (.I0(g1092),
        .I1(g1138),
        .I2(g1130),
        .I3(g1134),
        .I4(g1251),
        .I5(g1158),
        .O(g1149_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1149_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7525),
        .Q(g1149));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g114_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g114));
  LUT5 #(
    .INIT(32'hF8888888)) 
    g1153_i_1
       (.I0(g1077),
        .I1(g1084),
        .I2(g1158),
        .I3(g652),
        .I4(g1176),
        .O(g6856));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1153_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6856),
        .Q(g1153));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1153),
        .Q(g1154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1155_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1154),
        .Q(g1155));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1156_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1081),
        .Q(g1156));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1157_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1156),
        .Q(g1157));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1158_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1159),
        .Q(g1158));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1159_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1157),
        .Q(g1159));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1160_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1163),
        .Q(g1160));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1163_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1073),
        .Q(g1163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1166_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1167),
        .Q(g1166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1167_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1170),
        .Q(g1167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1170_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1173),
        .Q(g1170));
  LUT5 #(
    .INIT(32'h00000080)) 
    g1173_i_1
       (.I0(g1122),
        .I1(g1142),
        .I2(g1126),
        .I3(g1173_i_2_n_0),
        .I4(g1173_i_3_n_0),
        .O(g7217));
  LUT3 #(
    .INIT(8'h7F)) 
    g1173_i_2
       (.I0(g1118),
        .I1(g1110),
        .I2(g1114),
        .O(g1173_i_2_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1173_i_3
       (.I0(g1087),
        .I1(g1098),
        .I2(g1106),
        .I3(g1102),
        .O(g1173_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1173_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7217),
        .Q(g1173));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g1176_i_1
       (.I0(g1182),
        .I1(g1179),
        .I2(g1073),
        .I3(g1163),
        .I4(g1160),
        .I5(g1186),
        .O(g5172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1176_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5172),
        .Q(g1176));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1186),
        .Q(g1179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g117_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g114),
        .Q(g117));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1160),
        .Q(g1182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1155),
        .Q(g1185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1182),
        .Q(g1186));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1189_i_1
       (.I0(g1189_i_2_n_0),
        .I1(g1189_i_3_n_0),
        .I2(g1189_i_4_n_0),
        .I3(g1189_i_5_n_0),
        .O(g6392));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_2
       (.I0(g773),
        .I1(g1276),
        .I2(g771),
        .I3(g1284),
        .O(g1189_i_2_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1189_i_3
       (.I0(g770),
        .I1(g1288),
        .I2(g769),
        .I3(g1292),
        .O(g1189_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_4
       (.I0(g768),
        .I1(g1300),
        .I2(g1272),
        .I3(g774),
        .I4(g1280),
        .I5(g772),
        .O(g1189_i_4_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g1189_i_5
       (.I0(g1300),
        .I1(g768),
        .I2(g774),
        .I3(g1272),
        .I4(g767),
        .I5(g1296),
        .O(g1189_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1189_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6392),
        .Q(g1189));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g118_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g118));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1190_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .I3(g1357),
        .I4(g1360),
        .I5(g1190),
        .O(g8677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8677),
        .Q(g1190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1191_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g1191));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1192_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1191),
        .Q(g1192));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1193_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1192),
        .Q(g1193));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1194_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1193),
        .Q(g1194));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g1195));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1195),
        .Q(g1196));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1197_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1196),
        .Q(g1197));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1198_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1197),
        .Q(g1198));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g1199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g11_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g11),
        .Q(g11));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1199),
        .Q(g1200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1200),
        .Q(g1201));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1201),
        .Q(g1202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1203_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g1203));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1204_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1203),
        .Q(g1204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1204),
        .Q(g1205));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1206_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1205),
        .Q(g1206));
  LUT2 #(
    .INIT(4'hB)) 
    g1207_i_1
       (.I0(g1231),
        .I1(g1207),
        .O(g5173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5173),
        .Q(g1207));
  LUT3 #(
    .INIT(8'hBE)) 
    g1211_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .O(g5174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5174),
        .Q(g1211));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1214_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1211),
        .I3(g1207),
        .I4(g1214),
        .O(g5736));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5736),
        .Q(g1214));
  LUT5 #(
    .INIT(32'hBFFFEAAA)) 
    g1217_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1211),
        .I3(g1214),
        .I4(g1217),
        .O(g6377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1217_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6377),
        .Q(g1217));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g121_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g118),
        .Q(g121));
  LUT6 #(
    .INIT(64'hBFFFFFFFEAAAAAAA)) 
    g1220_i_1
       (.I0(g1231),
        .I1(g1214),
        .I2(g1211),
        .I3(g1207),
        .I4(g1217),
        .I5(g1220),
        .O(g6378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1220_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6378),
        .Q(g1220));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1223_i_1
       (.I0(g1231),
        .I1(g1217),
        .I2(g1207),
        .I3(g1223_i_2_n_0),
        .I4(g1220),
        .I5(g1223),
        .O(g6379));
  LUT2 #(
    .INIT(4'h7)) 
    g1223_i_2
       (.I0(g1214),
        .I1(g1211),
        .O(g1223_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1223_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6379),
        .Q(g1223));
  LUT3 #(
    .INIT(8'hBE)) 
    g1224_i_1
       (.I0(g1231),
        .I1(g1224_i_2_n_0),
        .I2(g1224),
        .O(g6857));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1224_i_2
       (.I0(g1223),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .I5(g1217),
        .O(g1224_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1224_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6857),
        .Q(g1224));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g1225_i_1
       (.I0(g1231),
        .I1(g1224),
        .I2(g1224_i_2_n_0),
        .I3(g1225),
        .O(g6858));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1225_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6858),
        .Q(g1225));
  LUT4 #(
    .INIT(16'hFBAE)) 
    g1226_i_1
       (.I0(g1231),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g6859));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    g1226_i_2
       (.I0(g1223),
        .I1(g1224),
        .I2(g1225),
        .I3(g1220),
        .I4(g1223_i_2_n_0),
        .I5(g1217),
        .O(g1226_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1226_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6859),
        .Q(g1226));
  LUT5 #(
    .INIT(32'hFBFFAEAA)) 
    g1227_i_1
       (.I0(g1231),
        .I1(g1226),
        .I2(g1226_i_2_n_0),
        .I3(g1207),
        .I4(g1227),
        .O(g7108));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1227_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7108),
        .Q(g1227));
  LUT6 #(
    .INIT(64'hFFBFFFFFAAEAAAAA)) 
    g1228_i_1
       (.I0(g1231),
        .I1(g1227),
        .I2(g1207),
        .I3(g1226_i_2_n_0),
        .I4(g1226),
        .I5(g1228),
        .O(g7109));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1228_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7109),
        .Q(g1228));
  LUT5 #(
    .INIT(32'h04444000)) 
    g1229_i_1
       (.I0(g1231),
        .I1(g1254),
        .I2(g1228),
        .I3(g1229_i_2_n_0),
        .I4(g1229),
        .O(g7110));
  LUT4 #(
    .INIT(16'h0800)) 
    g1229_i_2
       (.I0(g1227),
        .I1(g1207),
        .I2(g1226_i_2_n_0),
        .I3(g1226),
        .O(g1229_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1229_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7110),
        .Q(g1229));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g122_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g122));
  LUT4 #(
    .INIT(16'hEBAA)) 
    g1230_i_1
       (.I0(g1231),
        .I1(g1230),
        .I2(g1230_i_2_n_0),
        .I3(g1254),
        .O(g7300));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    g1230_i_2
       (.I0(g1226),
        .I1(g1226_i_2_n_0),
        .I2(g1229),
        .I3(g1227),
        .I4(g1228),
        .I5(g1207),
        .O(g1230_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1230_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7300),
        .Q(g1230));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1240_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1234),
        .Q(g1240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1243_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1240),
        .Q(g1243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1244_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1231),
        .Q(g1244));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1245_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1244),
        .Q(g1245));
  LUT2 #(
    .INIT(4'hB)) 
    g1247_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .O(g6380));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1247_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6380),
        .Q(g1247));
  LUT5 #(
    .INIT(32'hA0B0FFFF)) 
    g1250_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1263),
        .I2(g1247),
        .I3(g1257),
        .I4(g1253),
        .O(g7111));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1250_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7111),
        .Q(g1250));
  LUT4 #(
    .INIT(16'hCC04)) 
    g1251_i_1
       (.I0(g1257),
        .I1(g1247),
        .I2(g1263),
        .I3(g1254_i_2_n_0),
        .O(g6098));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1251_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6098),
        .Q(g1251));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1252_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1260),
        .Q(g1252));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1253_i_1
       (.I0(g1272),
        .I1(g1284),
        .I2(g1280),
        .I3(g1276),
        .I4(g1253_i_2_n_0),
        .O(g4681));
  LUT4 #(
    .INIT(16'h8000)) 
    g1253_i_2
       (.I0(g1296),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .O(g1253_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1253_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4681),
        .Q(g1253));
  LUT2 #(
    .INIT(4'hB)) 
    g1254_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1257),
        .O(g6381));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    g1254_i_2
       (.I0(g1226),
        .I1(g1228),
        .I2(g1223),
        .I3(g1230),
        .I4(g1254_i_3_n_0),
        .O(g1254_i_2_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1254_i_3
       (.I0(g1227),
        .I1(g1229),
        .I2(g1225),
        .I3(g1224),
        .O(g1254_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1254_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6381),
        .Q(g1254));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1257_i_1
       (.I0(g1217),
        .I1(g1220),
        .I2(g1214),
        .I3(g1211),
        .I4(g1207),
        .O(g5738));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1257_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5738),
        .Q(g1257));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g125_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g122),
        .Q(g125));
  LUT2 #(
    .INIT(4'hB)) 
    g1260_i_1
       (.I0(g1254_i_2_n_0),
        .I1(g1266),
        .O(g6382));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1260_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6382),
        .Q(g1260));
  LUT5 #(
    .INIT(32'h00008000)) 
    g1263_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5737));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1263_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5737),
        .Q(g1263));
  LUT5 #(
    .INIT(32'h00004000)) 
    g1266_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1220),
        .I3(g1217),
        .I4(g1207),
        .O(g5739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1266_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5739),
        .Q(g1266));
  LUT2 #(
    .INIT(4'h1)) 
    g1267_i_1
       (.I0(g1269),
        .I1(g1268),
        .O(g4656));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1267_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4656),
        .Q(g1267));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1268_i_1
       (.I0(g1227),
        .I1(g1230),
        .I2(g1224),
        .I3(g1228),
        .I4(g1268_i_2_n_0),
        .O(g5175));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1268_i_2
       (.I0(g1229),
        .I1(g1226),
        .I2(g1225),
        .I3(g1223),
        .O(g1268_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1268_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5175),
        .Q(g1268));
  LUT4 #(
    .INIT(16'hFFF7)) 
    g1269_i_1
       (.I0(g1211),
        .I1(g1214),
        .I2(g1217),
        .I3(g1220),
        .O(g5740));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1269_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5740),
        .Q(g1269));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g126_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g126));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1270_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1271),
        .Q(g1270));
  LUT2 #(
    .INIT(4'h2)) 
    g1271_i_1
       (.I0(g154),
        .I1(g1034),
        .O(g4792));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1271_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4792),
        .Q(g1271));
  LUT3 #(
    .INIT(8'h06)) 
    g1272_i_1
       (.I0(g1307),
        .I1(g1272),
        .I2(g1304),
        .O(g6383));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1272_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6383),
        .Q(g1272));
  LUT4 #(
    .INIT(16'h1540)) 
    g1276_i_1
       (.I0(g1304),
        .I1(g1272),
        .I2(g1307),
        .I3(g1276),
        .O(g6384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1276_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6384),
        .Q(g1276));
  LUT5 #(
    .INIT(32'h00007F80)) 
    g1280_i_1
       (.I0(g1276),
        .I1(g1307),
        .I2(g1272),
        .I3(g1280),
        .I4(g1304),
        .O(g7112));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1280_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7112),
        .Q(g1280));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1284_i_1
       (.I0(g1304),
        .I1(g1280),
        .I2(g1272),
        .I3(g1307),
        .I4(g1276),
        .I5(g1284),
        .O(g1284_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1284_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284_i_1_n_0),
        .Q(g1284));
  LUT6 #(
    .INIT(64'hFEBEBEBEBEBEBEBE)) 
    g1288_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1288_i_2_n_0),
        .I3(g1292),
        .I4(g1300),
        .I5(g1296),
        .O(g7527));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1288_i_2
       (.I0(g1307),
        .I1(g1272),
        .I2(g1284),
        .I3(g1280),
        .I4(g1276),
        .O(g1288_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1288_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7527),
        .Q(g1288));
  LUT3 #(
    .INIT(8'h41)) 
    g1292_i_1
       (.I0(g1304),
        .I1(g1300_i_2_n_0),
        .I2(g1292),
        .O(g7302));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7302),
        .Q(g1292));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    g1296_i_1
       (.I0(g1304),
        .I1(g1288),
        .I2(g1300),
        .I3(g1292),
        .I4(g1288_i_2_n_0),
        .I5(g1296),
        .O(g1296_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296_i_1_n_0),
        .Q(g1296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g129_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g126),
        .Q(g129));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g12_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7048),
        .Q(g12));
  LUT4 #(
    .INIT(16'h00D2)) 
    g1300_i_1
       (.I0(g1292),
        .I1(g1300_i_2_n_0),
        .I2(g1300),
        .I3(g1304),
        .O(g7303));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    g1300_i_2
       (.I0(g1288),
        .I1(g1276),
        .I2(g1280),
        .I3(g1284),
        .I4(g1272),
        .I5(g1307),
        .O(g1300_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1300_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7303),
        .Q(g1300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1304_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1312),
        .Q(g1304));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1307_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1307));
  LUT3 #(
    .INIT(8'hBA)) 
    g1308_i_1
       (.I0(g1236),
        .I1(g1034),
        .I2(g154),
        .O(g6385));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1308_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6385),
        .Q(g1308));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1309_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1308),
        .Q(g1309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g130_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g130));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1310_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1309),
        .Q(g1310));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1311_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1310),
        .Q(g1311));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1311),
        .Q(g1312));
  LUT3 #(
    .INIT(8'hA3)) 
    g1313_i_1
       (.I0(g145),
        .I1(g1313),
        .I2(g1329),
        .O(g5742));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5742),
        .Q(g1313));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1317_i_1
       (.I0(g141),
        .I1(g1329),
        .I2(g1317),
        .I3(g1313),
        .O(g5743));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5743),
        .Q(g1317));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1318_i_1
       (.I0(g137),
        .I1(g1329),
        .I2(g1318),
        .I3(g1317),
        .I4(g1313),
        .O(g6861));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1318_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6861),
        .Q(g1318));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1319_i_1
       (.I0(g133),
        .I1(g1329),
        .I2(g1319),
        .I3(g1318),
        .I4(g1317),
        .I5(g1313),
        .O(g7113));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1319_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7113),
        .Q(g1319));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1320_i_1
       (.I0(g129),
        .I1(g1329),
        .I2(g1320),
        .I3(g1320_i_2_n_0),
        .O(g7114));
  LUT4 #(
    .INIT(16'h8000)) 
    g1320_i_2
       (.I0(g1319),
        .I1(g1318),
        .I2(g1317),
        .I3(g1313),
        .O(g1320_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1320_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7114),
        .Q(g1320));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1321_i_1
       (.I0(g125),
        .I1(g1329),
        .I2(g1321),
        .I3(g1320_i_2_n_0),
        .I4(g1320),
        .O(g7115));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1321_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7115),
        .Q(g1321));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1322_i_1
       (.I0(g121),
        .I1(g1329),
        .I2(g1322),
        .I3(g1321),
        .I4(g1320),
        .I5(g1320_i_2_n_0),
        .O(g7116));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1322_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7116),
        .Q(g1322));
  LUT5 #(
    .INIT(32'hB88BB8B8)) 
    g1323_i_1
       (.I0(g117),
        .I1(g1329),
        .I2(g1323),
        .I3(g1323_i_2_n_0),
        .I4(g1320_i_2_n_0),
        .O(g7117));
  LUT3 #(
    .INIT(8'h7F)) 
    g1323_i_2
       (.I0(g1322),
        .I1(g1320),
        .I2(g1321),
        .O(g1323_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1323_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7117),
        .Q(g1323));
  LUT4 #(
    .INIT(16'h8BB8)) 
    g1324_i_1
       (.I0(g113),
        .I1(g1329),
        .I2(g1324),
        .I3(g1324_i_2_n_0),
        .O(g7118));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1324_i_2
       (.I0(g1320_i_2_n_0),
        .I1(g1323),
        .I2(g1322),
        .I3(g1320),
        .I4(g1321),
        .O(g1324_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1324_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7118),
        .Q(g1324));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1325_i_1
       (.I0(g108),
        .I1(g1329),
        .I2(g1325),
        .I3(g1324_i_2_n_0),
        .I4(g1324),
        .O(g7305));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1325_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7305),
        .Q(g1325));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1326_i_1
       (.I0(g103),
        .I1(g1329),
        .I2(g1326),
        .I3(g1324),
        .I4(g1324_i_2_n_0),
        .I5(g1325),
        .O(g7306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1326_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7306),
        .Q(g1326));
  LUT5 #(
    .INIT(32'h8BB8B8B8)) 
    g1327_i_1
       (.I0(g98),
        .I1(g1329),
        .I2(g1327),
        .I3(g1326),
        .I4(g1327_i_2_n_0),
        .O(g7307));
  LUT3 #(
    .INIT(8'h80)) 
    g1327_i_2
       (.I0(g1325),
        .I1(g1324_i_2_n_0),
        .I2(g1324),
        .O(g1327_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1327_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7307),
        .Q(g1327));
  LUT6 #(
    .INIT(64'h8BB8B8B8B8B8B8B8)) 
    g1328_i_1
       (.I0(g93),
        .I1(g1329),
        .I2(g1328),
        .I3(g1326),
        .I4(g1327),
        .I5(g1327_i_2_n_0),
        .O(g7309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1328_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7309),
        .Q(g1328));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1329_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1267),
        .Q(g1329));
  LUT2 #(
    .INIT(4'h2)) 
    g1330_i_1
       (.I0(g1247),
        .I1(g1330),
        .O(g6862));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1330_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6862),
        .Q(g1330));
  LUT3 #(
    .INIT(8'h60)) 
    g1333_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1247),
        .O(g1333_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1333_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1333_i_1_n_0),
        .Q(g1333));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1336_i_1
       (.I0(g1247),
        .I1(g1330),
        .I2(g1333),
        .I3(g1336),
        .O(g6864));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1336_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6864),
        .Q(g1336));
  LUT5 #(
    .INIT(32'h7F800000)) 
    g1339_i_1
       (.I0(g1333),
        .I1(g1330),
        .I2(g1336),
        .I3(g1339),
        .I4(g1247),
        .O(g1339_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1339_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1339_i_1_n_0),
        .Q(g1339));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g133_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g130),
        .Q(g133));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1342_i_1
       (.I0(g1247),
        .I1(g1339),
        .I2(g1336),
        .I3(g1330),
        .I4(g1333),
        .I5(g1342),
        .O(g7119));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1342_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7119),
        .Q(g1342));
  LUT4 #(
    .INIT(16'hA208)) 
    g1345_i_1
       (.I0(g1247),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1345),
        .O(g7528));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g1345_i_2
       (.I0(g1339),
        .I1(g1336),
        .I2(g1330),
        .I3(g1333),
        .O(g1345_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1345_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7528),
        .Q(g1345));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1348_i_1
       (.I0(g1247),
        .I1(g1345_i_2_n_0),
        .I2(g1342),
        .I3(g1345),
        .I4(g1348),
        .O(g7529));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1348_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7529),
        .Q(g1348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g134_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g134));
  LUT6 #(
    .INIT(64'hF7FF080000000000)) 
    g1351_i_1
       (.I0(g1345),
        .I1(g1342),
        .I2(g1345_i_2_n_0),
        .I3(g1348),
        .I4(g1351),
        .I5(g1247),
        .O(g1351_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1351_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1351_i_1_n_0),
        .Q(g1351));
  LUT3 #(
    .INIT(8'h28)) 
    g1354_i_1
       (.I0(g1247),
        .I1(g1354_i_2_n_0),
        .I2(g1354),
        .O(g7768));
  LUT5 #(
    .INIT(32'h00800000)) 
    g1354_i_2
       (.I0(g1342),
        .I1(g1348),
        .I2(g1351),
        .I3(g1345_i_2_n_0),
        .I4(g1345),
        .O(g1354_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7768),
        .Q(g1354));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1357_i_1
       (.I0(g1247),
        .I1(g1354),
        .I2(g1354_i_2_n_0),
        .I3(g1357),
        .O(g8675));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1357_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8675),
        .Q(g1357));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1360_i_1
       (.I0(g1247),
        .I1(g1357),
        .I2(g1354),
        .I3(g1354_i_2_n_0),
        .I4(g1360),
        .O(g8676));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1360_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8676),
        .Q(g1360));
  LUT2 #(
    .INIT(4'h6)) 
    g1363_i_1
       (.I0(g1227),
        .I1(g599),
        .O(g6877));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1363_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6877),
        .Q(g1363));
  LUT2 #(
    .INIT(4'h6)) 
    g1364_i_1
       (.I0(g1228),
        .I1(g598),
        .O(g6878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1364_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6878),
        .Q(g1364));
  LUT2 #(
    .INIT(4'h6)) 
    g1365_i_1
       (.I0(g1229),
        .I1(g597),
        .O(g6867));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1365_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6867),
        .Q(g1365));
  LUT2 #(
    .INIT(4'h6)) 
    g1366_i_1
       (.I0(g1230),
        .I1(g596),
        .O(g6866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1366_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6866),
        .Q(g1366));
  LUT2 #(
    .INIT(4'h6)) 
    g1367_i_1
       (.I0(g1223),
        .I1(g603),
        .O(g6873));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1367_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6873),
        .Q(g1367));
  LUT2 #(
    .INIT(4'h6)) 
    g1368_i_1
       (.I0(g1224),
        .I1(g602),
        .O(g6874));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6874),
        .Q(g1368));
  LUT2 #(
    .INIT(4'h6)) 
    g1369_i_1
       (.I0(g1225),
        .I1(g601),
        .O(g6875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1369_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6875),
        .Q(g1369));
  LUT2 #(
    .INIT(4'h6)) 
    g1370_i_1
       (.I0(g1226),
        .I1(g600),
        .O(g6876));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1370_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6876),
        .Q(g1370));
  LUT2 #(
    .INIT(4'h6)) 
    g1371_i_1
       (.I0(g1211),
        .I1(g607),
        .O(g6868));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6868),
        .Q(g1371));
  LUT2 #(
    .INIT(4'h6)) 
    g1372_i_1
       (.I0(g1214),
        .I1(g606),
        .O(g6870));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1372_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6870),
        .Q(g1372));
  LUT2 #(
    .INIT(4'h6)) 
    g1373_i_1
       (.I0(g1217),
        .I1(g605),
        .O(g6871));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6871),
        .Q(g1373));
  LUT2 #(
    .INIT(4'h6)) 
    g1374_i_1
       (.I0(g1220),
        .I1(g604),
        .O(g6872));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6872),
        .Q(g1374));
  LUT2 #(
    .INIT(4'h6)) 
    g1375_i_1
       (.I0(g1207),
        .I1(g608),
        .O(g6869));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6869),
        .Q(g1375));
  LUT2 #(
    .INIT(4'h6)) 
    g1376_i_1
       (.I0(g1227),
        .I1(g612),
        .O(g6890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6890),
        .Q(g1376));
  LUT2 #(
    .INIT(4'h6)) 
    g1377_i_1
       (.I0(g1228),
        .I1(g611),
        .O(g6891));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6891),
        .Q(g1377));
  LUT2 #(
    .INIT(4'h6)) 
    g1378_i_1
       (.I0(g1229),
        .I1(g610),
        .O(g6880));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1378_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6880),
        .Q(g1378));
  LUT2 #(
    .INIT(4'h6)) 
    g1379_i_1
       (.I0(g1230),
        .I1(g609),
        .O(g6879));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1379_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6879),
        .Q(g1379));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g137_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g134),
        .Q(g137));
  LUT2 #(
    .INIT(4'h6)) 
    g1380_i_1
       (.I0(g1223),
        .I1(g616),
        .O(g6886));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1380_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6886),
        .Q(g1380));
  LUT2 #(
    .INIT(4'h6)) 
    g1381_i_1
       (.I0(g1224),
        .I1(g615),
        .O(g6887));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1381_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6887),
        .Q(g1381));
  LUT2 #(
    .INIT(4'h6)) 
    g1382_i_1
       (.I0(g1225),
        .I1(g614),
        .O(g6888));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1382_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6888),
        .Q(g1382));
  LUT2 #(
    .INIT(4'h6)) 
    g1383_i_1
       (.I0(g1226),
        .I1(g613),
        .O(g6889));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1383_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6889),
        .Q(g1383));
  LUT2 #(
    .INIT(4'h6)) 
    g1384_i_1
       (.I0(g1211),
        .I1(g620),
        .O(g6881));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1384_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6881),
        .Q(g1384));
  LUT2 #(
    .INIT(4'h6)) 
    g1385_i_1
       (.I0(g1214),
        .I1(g619),
        .O(g6883));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1385_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6883),
        .Q(g1385));
  LUT2 #(
    .INIT(4'h6)) 
    g1386_i_1
       (.I0(g1217),
        .I1(g618),
        .O(g6884));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1386_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6884),
        .Q(g1386));
  LUT2 #(
    .INIT(4'h6)) 
    g1387_i_1
       (.I0(g1220),
        .I1(g617),
        .O(g6885));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1387_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6885),
        .Q(g1387));
  LUT2 #(
    .INIT(4'h6)) 
    g1388_i_1
       (.I0(g1207),
        .I1(g621),
        .O(g6882));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1388_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6882),
        .Q(g1388));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g1389_i_1
       (.I0(g1389_i_2_n_0),
        .I1(g2262),
        .I2(g1378),
        .I3(g1377),
        .I4(g1376),
        .I5(g1379),
        .O(g4658));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g1389_i_2
       (.I0(g1383),
        .I1(g1380),
        .I2(g1381),
        .I3(g1382),
        .I4(g1388),
        .O(g1389_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g1389_i_3
       (.I0(g1386),
        .I1(g1385),
        .I2(g1384),
        .I3(g1387),
        .O(g2262));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1389_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4658),
        .Q(g1389));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g138_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g138));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1390_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1251),
        .Q(g1390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1391_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1390),
        .Q(g1391));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1392_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g1392));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g16),
        .Q(g1393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g1394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1393),
        .Q(g1395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1250),
        .Q(g1396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g1397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1396),
        .Q(g1398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1399_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7731),
        .Q(g1399));
  LUT4 #(
    .INIT(16'h00F2)) 
    g13_i_1
       (.I0(g1324_i_2_n_0),
        .I1(g13_i_2_n_0),
        .I2(g13),
        .I3(g1329),
        .O(g7308));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    g13_i_2
       (.I0(g1328),
        .I1(g1327),
        .I2(g1326),
        .I3(g1324),
        .I4(g1325),
        .O(g13_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g13_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7308),
        .Q(g13));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1400_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g1400));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1401_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1399),
        .Q(g1401));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g1402_i_1
       (.I0(g1402_i_2_n_0),
        .I1(g763),
        .I2(g1345),
        .I3(g762),
        .I4(g1348),
        .I5(g1402_i_3_n_0),
        .O(g6391));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_2
       (.I0(g765),
        .I1(g1339),
        .I2(g764),
        .I3(g1342),
        .O(g1402_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF6)) 
    g1402_i_3
       (.I0(g1336),
        .I1(g766),
        .I2(g1330),
        .I3(g1333),
        .I4(g1402_i_4_n_0),
        .I5(g1402_i_5_n_0),
        .O(g1402_i_3_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_4
       (.I0(g761),
        .I1(g1351),
        .I2(g759),
        .I3(g1357),
        .O(g1402_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g1402_i_5
       (.I0(g760),
        .I1(g1354),
        .I2(g758),
        .I3(g1360),
        .O(g1402_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1402_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6391),
        .Q(g1402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1403_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1402),
        .Q(g1403));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1404_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1403),
        .Q(g1404));
  LUT4 #(
    .INIT(16'h0007)) 
    g1405_i_1
       (.I0(g1408),
        .I1(g1405),
        .I2(g1428),
        .I3(g1429),
        .O(g5744));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1405_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5744),
        .Q(g1405));
  LUT3 #(
    .INIT(8'hFE)) 
    g1408_i_1
       (.I0(g1405),
        .I1(g1428),
        .I2(g1429),
        .O(g5177));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1408_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5177),
        .Q(g1408));
  LUT4 #(
    .INIT(16'h8BBB)) 
    g1409_i_1
       (.I0(g1409),
        .I1(g1416),
        .I2(g1412),
        .I3(g1405),
        .O(g5178));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1409_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5178),
        .Q(g1409));
  LUT4 #(
    .INIT(16'h0111)) 
    g1412_i_1
       (.I0(g1430),
        .I1(g1431),
        .I2(g1415),
        .I3(g1412),
        .O(g5745));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1412_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5745),
        .Q(g1412));
  LUT3 #(
    .INIT(8'hFE)) 
    g1415_i_1
       (.I0(g1412),
        .I1(g1430),
        .I2(g1431),
        .O(g5180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1415_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5180),
        .Q(g1415));
  LUT3 #(
    .INIT(8'hF1)) 
    g1416_i_1
       (.I0(g1421),
        .I1(g1416),
        .I2(g1424),
        .O(g4665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1416_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4665),
        .Q(g1416));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g141_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g138),
        .Q(g141));
  LUT3 #(
    .INIT(8'h02)) 
    g1421_i_1
       (.I0(g1416),
        .I1(g1421),
        .I2(g1424),
        .O(g1421_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1421_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1421_i_1_n_0),
        .Q(g1421));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1424_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1424));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1428_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1424),
        .Q(g1428));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1429_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1236),
        .Q(g1429));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g142_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g142));
  LUT1 #(
    .INIT(2'h1)) 
    g1430_i_1
       (.I0(g1252),
        .O(g4666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1430_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1430));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1431_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1243),
        .Q(g1431));
  LUT4 #(
    .INIT(16'h0038)) 
    g1432_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1432_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5183),
        .Q(g1432));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1435_i_1
       (.I0(g1439),
        .I1(g1432),
        .I2(g1443),
        .I3(g1435),
        .O(g1435_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1435_i_1_n_0),
        .Q(g1435));
  LUT4 #(
    .INIT(16'h0026)) 
    g1439_i_1
       (.I0(g1435),
        .I1(g1439),
        .I2(g1432),
        .I3(g1443),
        .O(g5182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1439_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5182),
        .Q(g1439));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1443_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4666),
        .Q(g1443));
  LUT4 #(
    .INIT(16'hF8FF)) 
    g1444_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1459),
        .I3(g1444),
        .O(g1444_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1444_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1444_i_1_n_0),
        .Q(g1444));
  LUT4 #(
    .INIT(16'h0026)) 
    g1450_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5186));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1450_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5186),
        .Q(g1450));
  LUT4 #(
    .INIT(16'h0038)) 
    g1454_i_1
       (.I0(g1444),
        .I1(g1450),
        .I2(g1454),
        .I3(g1459),
        .O(g5187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5187),
        .Q(g1454));
  LUT1 #(
    .INIT(2'h1)) 
    g1459_i_1
       (.I0(g1260),
        .O(g3863));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1459_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3863),
        .Q(g1459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g145_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g142),
        .Q(g145));
  LUT3 #(
    .INIT(8'h02)) 
    g1460_i_1
       (.I0(g1450),
        .I1(g1454),
        .I2(g1444),
        .O(g4668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1460_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4668),
        .Q(g1460));
  LUT3 #(
    .INIT(8'h08)) 
    g1461_i_1
       (.I0(g1454),
        .I1(g1444),
        .I2(g1450),
        .O(g1461_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1461_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1461_i_1_n_0),
        .Q(g1461));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g1462_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .I5(g1462),
        .O(g8678));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1462_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8678),
        .Q(g1462));
  LUT3 #(
    .INIT(8'h28)) 
    g1467_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1467_i_2_n_0),
        .I2(g1467),
        .O(g8875));
  LUT5 #(
    .INIT(32'h80000000)) 
    g1467_i_2
       (.I0(g1462),
        .I1(g1519),
        .I2(g1514),
        .I3(g1509),
        .I4(g1509_i_2_n_0),
        .O(g1467_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1467_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8875),
        .Q(g1467));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g146_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g146));
  LUT3 #(
    .INIT(8'h28)) 
    g1472_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1472_i_2_n_0),
        .O(g8960));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g1472_i_2
       (.I0(g1467),
        .I1(g1514),
        .I2(g1509_i_2_n_0),
        .I3(g1509),
        .I4(g1519),
        .I5(g1462),
        .O(g1472_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1472_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8960),
        .Q(g1472));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1477_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1472),
        .I2(g1467),
        .I3(g1467_i_2_n_0),
        .I4(g1477),
        .O(g9036));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9036),
        .Q(g1477));
  LUT3 #(
    .INIT(8'h82)) 
    g1481_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .O(g7769));
  LUT5 #(
    .INIT(32'h0000FF9F)) 
    g1481_i_2
       (.I0(g1524),
        .I1(g1513),
        .I2(g150),
        .I3(g1034),
        .I4(g1486_i_2_n_0),
        .O(g1481_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1481_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7769),
        .Q(g1481));
  LUT5 #(
    .INIT(32'h3C3C553C)) 
    g1486_i_1
       (.I0(g1524),
        .I1(g1486),
        .I2(g1486_i_2_n_0),
        .I3(g150),
        .I4(g1034),
        .O(g8226));
  LUT6 #(
    .INIT(64'h0202000200020002)) 
    g1486_i_2
       (.I0(g1486_i_3_n_0),
        .I1(g1486_i_4_n_0),
        .I2(g1486_i_5_n_0),
        .I3(g174),
        .I4(g1477),
        .I5(g1504),
        .O(g1486_i_2_n_0));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    g1486_i_3
       (.I0(g174),
        .I1(g1514),
        .I2(g1481),
        .I3(g1489),
        .I4(g150),
        .I5(g1034),
        .O(g1486_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g1486_i_4
       (.I0(g1472),
        .I1(g1462),
        .I2(g1499),
        .O(g1486_i_4_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g1486_i_5
       (.I0(g1519),
        .I1(g1251),
        .I2(g1467),
        .I3(g1494),
        .O(g1486_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1486_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8226),
        .Q(g1486));
  LUT4 #(
    .INIT(16'hA208)) 
    g1489_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1481),
        .I2(g1251),
        .I3(g1489),
        .O(g7770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1489_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7770),
        .Q(g1489));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1494_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1251),
        .I2(g1481),
        .I3(g1489),
        .I4(g1494),
        .O(g7771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1494_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7771),
        .Q(g1494));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    g1499_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1489),
        .I2(g1481),
        .I3(g1251),
        .I4(g1494),
        .I5(g1499),
        .O(g7772));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1499_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7772),
        .Q(g1499));
  LUT3 #(
    .INIT(8'h28)) 
    g1504_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1504_i_2_n_0),
        .I2(g1504),
        .O(g7773));
  LUT5 #(
    .INIT(32'h40000000)) 
    g1504_i_2
       (.I0(g1251),
        .I1(g1499),
        .I2(g1489),
        .I3(g1481),
        .I4(g1494),
        .O(g1504_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1504_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7773),
        .Q(g1504));
  LUT3 #(
    .INIT(8'h28)) 
    g1509_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .O(g7774));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    g1509_i_2
       (.I0(g1494),
        .I1(g1481),
        .I2(g1489),
        .I3(g1499),
        .I4(g1251),
        .I5(g1504),
        .O(g1509_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1509_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7774),
        .Q(g1509));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g150_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g150));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1513_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1524),
        .Q(g1513));
  LUT4 #(
    .INIT(16'h2A80)) 
    g1514_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509_i_2_n_0),
        .I2(g1509),
        .I3(g1514),
        .O(g7775));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1514_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7775),
        .Q(g1514));
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    g1519_i_1
       (.I0(g1481_i_2_n_0),
        .I1(g1509),
        .I2(g1509_i_2_n_0),
        .I3(g1514),
        .I4(g1519),
        .O(g8227));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1519_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8227),
        .Q(g1519));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1524_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g1524));
  LUT4 #(
    .INIT(16'hA208)) 
    g1528_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1532),
        .I2(g1251),
        .I3(g1528),
        .O(g7776));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1528_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7776),
        .Q(g1528));
  LUT3 #(
    .INIT(8'h82)) 
    g1532_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .O(g7781));
  LUT3 #(
    .INIT(8'h15)) 
    g1532_i_2
       (.I0(g1553),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g1532_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1532_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7781),
        .Q(g1532));
  LUT5 #(
    .INIT(32'h8AAA2000)) 
    g1537_i_1
       (.I0(g1532_i_2_n_0),
        .I1(g1251),
        .I2(g1532),
        .I3(g1528),
        .I4(g1537),
        .O(g7777));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1537_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7777),
        .Q(g1537));
  LUT6 #(
    .INIT(64'hF7FF0800FFFFFFFF)) 
    g1541_i_1
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1532_i_2_n_0),
        .O(g7778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1541_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7778),
        .Q(g1541));
  LUT4 #(
    .INIT(16'hEFFC)) 
    g1545_i_1
       (.I0(g1549),
        .I1(g1553),
        .I2(g1545_i_2_n_0),
        .I3(g1545),
        .O(g7779));
  LUT5 #(
    .INIT(32'h08000000)) 
    g1545_i_2
       (.I0(g1541),
        .I1(g1537),
        .I2(g1251),
        .I3(g1532),
        .I4(g1528),
        .O(g1545_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1545_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7779),
        .Q(g1545));
  LUT3 #(
    .INIT(8'h14)) 
    g1549_i_1
       (.I0(g1553),
        .I1(g1549_i_2_n_0),
        .I2(g1549),
        .O(g7780));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    g1549_i_2
       (.I0(g1528),
        .I1(g1532),
        .I2(g1251),
        .I3(g1537),
        .I4(g1541),
        .I5(g1545),
        .O(g1549_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1549_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7780),
        .Q(g1549));
  LUT4 #(
    .INIT(16'h00E2)) 
    g154_i_1
       (.I0(g154),
        .I1(g162_i_1_n_0),
        .I2(g4),
        .I3(g172),
        .O(g7739));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g154_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7739),
        .Q(g154));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g158_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g158));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    g162_i_1
       (.I0(g58),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g162_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g162_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g162));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g168_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g16_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1404),
        .Q(g16));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g172_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1270),
        .Q(g172));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g173_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g173));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g174_reg
       (.C(blif_clk_net),
        .CE(g162_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g174));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g179_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g196),
        .Q(g179));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g180_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g187),
        .Q(g180));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g181_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g202),
        .Q(g181));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g182_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g207),
        .Q(g182));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g183_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g10),
        .Q(g183));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g184_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g185_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1034),
        .Q(g185));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g186_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g186));
  LUT4 #(
    .INIT(16'hF600)) 
    g187_i_1
       (.I0(g186),
        .I1(g1198),
        .I2(g187),
        .I3(g190),
        .O(g5730));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g187_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5730),
        .Q(g187));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g190_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g201),
        .Q(g190));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g195_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g195));
  LUT4 #(
    .INIT(16'hF600)) 
    g196_i_1
       (.I0(g195),
        .I1(g1194),
        .I2(g196),
        .I3(g190),
        .O(g5731));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g196_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5731),
        .Q(g196));
  LUT1 #(
    .INIT(2'h1)) 
    g199_i_1
       (.I0(g158),
        .O(g3832));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g199_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3832),
        .Q(g199));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g1_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1),
        .Q(g1));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g200_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g199),
        .Q(g200));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g201_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g200),
        .Q(g201));
  LUT4 #(
    .INIT(16'hF600)) 
    g202_i_1
       (.I0(g205),
        .I1(g1202),
        .I2(g202),
        .I3(g190),
        .O(g5732));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g202_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5732),
        .Q(g202));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g205_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g205));
  LUT4 #(
    .INIT(16'hF600)) 
    g207_i_1
       (.I0(g210),
        .I1(g1206),
        .I2(g207),
        .I3(g190),
        .O(g5733));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g207_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5733),
        .Q(g207));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    g20_i_1
       (.I0(g20_i_2_n_0),
        .I1(g627),
        .I2(g1345),
        .I3(g626),
        .I4(g1348),
        .I5(g20_i_3_n_0),
        .O(g6386));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_2
       (.I0(g629),
        .I1(g1339),
        .I2(g628),
        .I3(g1342),
        .O(g20_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFEFFFFFFFFEFFE)) 
    g20_i_3
       (.I0(g20_i_4_n_0),
        .I1(g20_i_5_n_0),
        .I2(g623),
        .I3(g1357),
        .I4(g622),
        .I5(g1360),
        .O(g20_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    g20_i_4
       (.I0(g631),
        .I1(g1333),
        .I2(g1336),
        .I3(g630),
        .I4(g1330),
        .I5(g632),
        .O(g20_i_4_n_0));
  LUT4 #(
    .INIT(16'h6FF6)) 
    g20_i_5
       (.I0(g624),
        .I1(g1354),
        .I2(g625),
        .I3(g1351),
        .O(g20_i_5_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g20_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6386),
        .Q(g20));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g210_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g210));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g211_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g211));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g212_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g212));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g213_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g213));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g214_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g214));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g215_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g215));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g216_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g211),
        .Q(g216));
  LUT2 #(
    .INIT(4'h2)) 
    g219_i_1
       (.I0(g290),
        .I1(g287),
        .O(g219_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g219_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g212),
        .Q(g219));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g21_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g21),
        .Q(g21));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g222_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g213),
        .Q(g222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g225_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g214),
        .Q(g225));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g228_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g215),
        .Q(g228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g22_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g22),
        .Q(g22));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g231_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g231));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g232_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g232));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g233_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g233));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g234_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g234));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g235_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g235));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g236_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g236));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g237_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g231),
        .Q(g237));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g23_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g23),
        .Q(g23));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g240_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g232),
        .Q(g240));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g243_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g233),
        .Q(g243));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g246_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g234),
        .Q(g246));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g249_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g235),
        .Q(g249));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g24_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g24),
        .Q(g24));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g252_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g236),
        .Q(g252));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g255_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g237),
        .Q(g255));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g258_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g240),
        .Q(g258));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g25_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g25),
        .Q(g25));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g261_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g243),
        .Q(g261));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g264_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g246),
        .Q(g264));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    g267_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g267_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g267_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g249),
        .Q(g267));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g26_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g26),
        .Q(g26));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g270_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g252),
        .Q(g270));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g273_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g273));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g274_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g274));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g275_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g273),
        .Q(g275));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g278_reg
       (.C(blif_clk_net),
        .CE(g219_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g274),
        .Q(g278));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g27_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g27),
        .Q(g27));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g281_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g275),
        .Q(g281));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g284_reg
       (.C(blif_clk_net),
        .CE(g267_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g278),
        .Q(g284));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g287_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1194),
        .Q(g287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g28_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g28),
        .Q(g28));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g290_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g287),
        .Q(g290));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g292_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g292));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g293_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g293));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g294_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g294));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g295_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g295));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g296_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g296));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g297_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g292),
        .Q(g297));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g29_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g29),
        .Q(g29));
  LUT6 #(
    .INIT(64'h5155515551550000)) 
    g2_i_1
       (.I0(g9299_INST_0_i_5_n_0),
        .I1(g9299_INST_0_i_4_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_2_n_0),
        .I4(g2_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9361));
  LUT6 #(
    .INIT(64'hFFFFEFEEFFFFFFFF)) 
    g2_i_2
       (.I0(g2_i_3_n_0),
        .I1(g9299_INST_0_i_8_n_0),
        .I2(g9305_INST_0_i_23_n_0),
        .I3(g222),
        .I4(g2_i_4_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g2_i_3
       (.I0(g9299_INST_0_i_30_n_0),
        .I1(g2_i_5_n_0),
        .I2(g2_i_6_n_0),
        .I3(g2_i_7_n_0),
        .I4(g611),
        .I5(g9299_INST_0_i_26_n_0),
        .O(g2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g2_i_4
       (.I0(g619),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g270),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_23_n_0),
        .O(g2_i_4_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_5
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g351),
        .I2(g706_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g134),
        .O(g2_i_5_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g2_i_6
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g573_i_2_n_0),
        .I4(g158),
        .O(g2_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    g2_i_7
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g68),
        .O(g2_i_7_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g2_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9361),
        .Q(g2));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g300_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g293),
        .Q(g300));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g303_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g294),
        .Q(g303));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g306_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g295),
        .Q(g306));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g309_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g296),
        .Q(g309));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g30_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g30),
        .Q(g30));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g312_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g312));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g313_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g313));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g314_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g314));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g315_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g315));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g316_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g316));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g317_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g317));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g318_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g312),
        .Q(g318));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g31_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g31),
        .Q(g31));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g321_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g313),
        .Q(g321));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g324_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g314),
        .Q(g324));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g327_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g315),
        .Q(g327));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g32_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g32),
        .Q(g32));
  LUT2 #(
    .INIT(4'h2)) 
    g330_i_1
       (.I0(g371),
        .I1(g368),
        .O(g330_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g330_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g316),
        .Q(g330));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g333_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g317),
        .Q(g333));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g336_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g318),
        .Q(g336));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g339_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g321),
        .Q(g339));
  LUT4 #(
    .INIT(16'hBFEA)) 
    g33_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .O(g5184));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g33_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5184),
        .Q(g33));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g342_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g324),
        .Q(g342));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g345_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g327),
        .Q(g345));
  LUT5 #(
    .INIT(32'h00100000)) 
    g348_i_1
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g348_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g348_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g330),
        .Q(g348));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g351_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g333),
        .Q(g351));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g354_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g354));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g355_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g355));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g356_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g354),
        .Q(g356));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g359_reg
       (.C(blif_clk_net),
        .CE(g330_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g355),
        .Q(g359));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g362_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g356),
        .Q(g362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g365_reg
       (.C(blif_clk_net),
        .CE(g348_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g359),
        .Q(g365));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g368_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1198),
        .Q(g368));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g371_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g368),
        .Q(g371));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g373_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g374_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g374));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g375_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g375));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g376_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g376));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g377_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g377));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g378_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g373),
        .Q(g378));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g37_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g37),
        .Q(g37));
  LUT2 #(
    .INIT(4'h2)) 
    g381_i_1
       (.I0(g452),
        .I1(g449),
        .O(g381_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g381_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g374),
        .Q(g381));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g384_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g375),
        .Q(g384));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g387_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g376),
        .Q(g387));
  LUT5 #(
    .INIT(32'hFFBFAAEA)) 
    g38_i_1
       (.I0(g1443),
        .I1(g1439),
        .I2(g1432),
        .I3(g33),
        .I4(g38),
        .O(g5746));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g38_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5746),
        .Q(g38));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g390_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g377),
        .Q(g390));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g393_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g393));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g394_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g394));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g395_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g395));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g396_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g396));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g397_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g397));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g398_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g398));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g399_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g393),
        .Q(g399));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g3_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9360),
        .Q(g3));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g402_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g394),
        .Q(g402));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g405_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g395),
        .Q(g405));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g408_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g396),
        .Q(g408));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g411_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g397),
        .Q(g411));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g414_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g398),
        .Q(g414));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g417_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g399),
        .Q(g417));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g41_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g41),
        .Q(g41));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g420_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g402),
        .Q(g420));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g423_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g405),
        .Q(g423));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g426_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g408),
        .Q(g426));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g429_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g411),
        .Q(g429));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g42_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g42),
        .Q(g42));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g432_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g414),
        .Q(g432));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g435_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g435));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g436_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g436));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g437_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g435),
        .Q(g437));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g440_reg
       (.C(blif_clk_net),
        .CE(g381_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g436),
        .Q(g440));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g443_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g437),
        .Q(g443));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g446_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g440),
        .Q(g446));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g449_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g449));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g44_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g44),
        .Q(g44));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g452_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g449),
        .Q(g452));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g454_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1230),
        .Q(g454));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g455_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1229),
        .Q(g455));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g456_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1228),
        .Q(g456));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g457_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1227),
        .Q(g457));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g458_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1226),
        .Q(g458));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g459_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g454),
        .Q(g459));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g45_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g45));
  LUT2 #(
    .INIT(4'h2)) 
    g462_i_1
       (.I0(g533),
        .I1(g530),
        .O(g462_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g462_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g455),
        .Q(g462));
  LUT2 #(
    .INIT(4'h6)) 
    g4655_INST_0
       (.I0(g940),
        .I1(g936),
        .O(g4655));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g4657_INST_0
       (.I0(g4657_INST_0_i_1_n_0),
        .I1(g2206),
        .I2(g1374),
        .I3(g1372),
        .I4(g1371),
        .I5(g1373),
        .O(g4657));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g4657_INST_0_i_1
       (.I0(g1370),
        .I1(g1367),
        .I2(g1368),
        .I3(g1369),
        .I4(g1375),
        .O(g4657_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g4657_INST_0_i_2
       (.I0(g1366),
        .I1(g1364),
        .I2(g1363),
        .I3(g1365),
        .O(g2206));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g465_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g456),
        .Q(g465));
  LUT2 #(
    .INIT(4'h2)) 
    g4660_INST_0
       (.I0(g1392),
        .I1(g1391),
        .O(g4660));
  LUT2 #(
    .INIT(4'h2)) 
    g4661_INST_0
       (.I0(g1394),
        .I1(g1395),
        .O(g4661));
  LUT2 #(
    .INIT(4'h2)) 
    g4663_INST_0
       (.I0(g1397),
        .I1(g1398),
        .O(g4663));
  LUT2 #(
    .INIT(4'h2)) 
    g4664_INST_0
       (.I0(g1400),
        .I1(g1401),
        .O(g4664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g468_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g457),
        .Q(g468));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g46_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g45),
        .Q(g46));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g471_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g458),
        .Q(g471));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g474_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1225),
        .Q(g474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g475_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1224),
        .Q(g475));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g476_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1223),
        .Q(g476));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g477_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1220),
        .Q(g477));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g478_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1217),
        .Q(g478));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g479_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1214),
        .Q(g479));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    g47_i_1
       (.I0(g9378_INST_0_i_4_n_0),
        .I1(g47_i_2_n_0),
        .I2(g47_i_3_n_0),
        .I3(g9378_INST_0_i_2_n_0),
        .I4(g44),
        .I5(g7480),
        .O(g9389));
  LUT6 #(
    .INIT(64'hFFFFFFF044444444)) 
    g47_i_2
       (.I0(g9378_INST_0_i_8_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g47_i_4_n_0),
        .I4(g47_i_5_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000FF10FF10)) 
    g47_i_3
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_3_n_0),
        .I2(g9378_INST_0_i_24_n_0),
        .I3(g9299_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g47_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    g47_i_4
       (.I0(g47_i_6_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_26_n_0),
        .I3(g9378_INST_0_i_12_n_0),
        .I4(g9378_INST_0_i_13_n_0),
        .O(g47_i_4_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g47_i_5
       (.I0(g9378_INST_0_i_14_n_0),
        .I1(g47_i_7_n_0),
        .I2(g9297_INST_0_i_11_n_0),
        .I3(g573),
        .I4(g9378_INST_0_i_32_n_0),
        .I5(g429),
        .O(g47_i_5_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g47_i_6
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g348),
        .I2(g180),
        .I3(g9310_INST_0_i_14_n_0),
        .I4(g267),
        .I5(g9299_INST_0_i_24_n_0),
        .O(g47_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g47_i_7
       (.I0(g9305_INST_0_i_23_n_0),
        .I1(g219),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g597),
        .O(g47_i_7_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g47_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9389),
        .Q(g47));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g480_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g474),
        .Q(g480));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g483_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g475),
        .Q(g483));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g486_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g476),
        .Q(g486));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g489_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g477),
        .Q(g489));
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g48_i_1
       (.I0(g9280_INST_0_i_1_n_0),
        .O(g9362));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g48_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9362),
        .Q(g48));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g492_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g478),
        .Q(g492));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g495_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g479),
        .Q(g495));
  LUT5 #(
    .INIT(32'h00001000)) 
    g498_i_1
       (.I0(g498_i_2_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .O(g498_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    g498_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g52),
        .O(g498_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g498_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g480),
        .Q(g498));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    g4_i_1
       (.I0(g9305_INST_0_i_5_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g4_i_2_n_0),
        .I3(g9305_INST_0_i_12_n_0),
        .I4(g9305_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_1_n_0),
        .O(g9372));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g4_i_2
       (.I0(g9305_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_15_n_0),
        .I2(g618),
        .I3(g4_i_3_n_0),
        .I4(g95),
        .I5(g9305_INST_0_i_13_n_0),
        .O(g4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g4_i_3
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g4_i_3_n_0));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g4_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9372),
        .Q(g4));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g501_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g483),
        .Q(g501));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g504_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g486),
        .Q(g504));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g507_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g489),
        .Q(g507));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g510_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g492),
        .Q(g510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g513_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g495),
        .Q(g513));
  LUT3 #(
    .INIT(8'h80)) 
    g5164_INST_0
       (.I0(g889),
        .I1(g887),
        .I2(g888),
        .O(g5164));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g516_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1211),
        .Q(g516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g517_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1207),
        .Q(g517));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g518_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g516),
        .Q(g518));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g521_reg
       (.C(blif_clk_net),
        .CE(g462_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g517),
        .Q(g521));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g524_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g518),
        .Q(g524));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g527_reg
       (.C(blif_clk_net),
        .CE(g498_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g521),
        .Q(g527));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g52_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g52));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g530_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1202),
        .Q(g530));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g533_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g530),
        .Q(g533));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g535_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1280),
        .Q(g535));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g536_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g535),
        .Q(g536));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g539_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1276),
        .Q(g539));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g540_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g539),
        .Q(g540));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g543_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1272),
        .Q(g543));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g544_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g543),
        .Q(g544));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g547_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g536),
        .Q(g547));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g550_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g540),
        .Q(g550));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g553_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g544),
        .Q(g553));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g556_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1296),
        .Q(g556));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g557_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g556),
        .Q(g557));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g55_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7480),
        .Q(g55));
  LUT2 #(
    .INIT(4'h2)) 
    g560_i_1
       (.I0(g595),
        .I1(g576),
        .O(g560_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g560_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g587),
        .Q(g560));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g563_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g557),
        .Q(g563));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g566_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1300),
        .Q(g566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g567_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g566),
        .Q(g567));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g570_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g567),
        .Q(g570));
  LUT5 #(
    .INIT(32'h00000004)) 
    g573_i_1
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g573_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g573_i_2
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g86),
        .I2(g83),
        .I3(g52),
        .I4(g80),
        .O(g573_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g573_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g560),
        .Q(g573));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g576_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1206),
        .Q(g576));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g579_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1292),
        .Q(g579));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g580_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g579),
        .Q(g580));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g583_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1288),
        .Q(g583));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g584_reg
       (.C(blif_clk_net),
        .CE(g560_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g583),
        .Q(g584));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g587_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1284),
        .Q(g587));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g588_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g580),
        .Q(g588));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g58_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(1'b0),
        .Q(g58));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g591_reg
       (.C(blif_clk_net),
        .CE(g573_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g584),
        .Q(g591));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g595_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g576),
        .Q(g595));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g596_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g596));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g597_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g597));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g598_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g599_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g599));
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT1 #(
    .INIT(2'h1)) 
    g5_i_1
       (.I0(g9308_INST_0_i_1_n_0),
        .O(g9373));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g5_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9373),
        .Q(g5));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g600_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g600));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g601_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g601));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g602_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g602));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g603_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g603));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g604_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g604));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g605_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g605));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g606_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g606));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g607_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g607));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g608_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g608));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g609_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g609));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g610_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g610));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g611_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g611));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g612_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g612));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g613_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g613));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g614_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g614));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g615_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g615));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g616_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g616));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g617_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g617));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g618_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g618));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g619_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g619));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g620_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g620));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g621_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g621));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g622_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g622));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g623_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g623));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g624_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g624));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g625_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g625));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g626_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g626));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g627_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g627));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g628_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g628));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g629_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g629));
  LUT5 #(
    .INIT(32'h00000004)) 
    g62_i_1
       (.I0(g55),
        .I1(g44),
        .I2(g45),
        .I3(g42),
        .I4(g41),
        .O(g7367));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g62_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7367),
        .Q(g62));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g630_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g630));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g631_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g631));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g632_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g632));
  LUT1 #(
    .INIT(2'h1)) 
    g646_i_1
       (.I0(g1158),
        .O(g4652));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g646_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4652),
        .Q(g646));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g652_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g646),
        .Q(g652));
  LUT2 #(
    .INIT(4'hE)) 
    g65_i_1
       (.I0(g58),
        .I1(g65),
        .O(g4598));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g65_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4598),
        .Q(g65));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g661_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g661));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g665_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g669_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g673_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g673));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g677_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g677));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g681_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g681));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g6849_INST_0
       (.I0(g6849_INST_0_i_1_n_0),
        .I1(g6849_INST_0_i_2_n_0),
        .I2(g6849_INST_0_i_3_n_0),
        .I3(g6849_INST_0_i_4_n_0),
        .I4(g6849_INST_0_i_5_n_0),
        .I5(g778),
        .O(g6849));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_1
       (.I0(g896),
        .I1(g834),
        .I2(g921),
        .I3(g849),
        .I4(g891),
        .I5(g831),
        .O(g6849_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_2
       (.I0(g849),
        .I1(g921),
        .I2(g837),
        .I3(g901),
        .I4(g911),
        .I5(g843),
        .O(g6849_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_3
       (.I0(g846),
        .I1(g916),
        .I2(g901),
        .I3(g837),
        .I4(g883),
        .I5(g852),
        .O(g6849_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFFFFFF22F2)) 
    g6849_INST_0_i_4
       (.I0(g916),
        .I1(g846),
        .I2(g834),
        .I3(g896),
        .I4(g840),
        .I5(g906),
        .O(g6849_INST_0_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g6849_INST_0_i_5
       (.I0(g887),
        .I1(g889),
        .I2(g888),
        .O(g6849_INST_0_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g6850_INST_0
       (.I0(g43),
        .O(g6850));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g685_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g685));
  LUT1 #(
    .INIT(2'h1)) 
    g6895_INST_0
       (.I0(g689),
        .O(g6895));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    g689_i_1
       (.I0(g689_i_2_n_0),
        .I1(g648),
        .I2(g685),
        .I3(g702),
        .I4(g718),
        .I5(g689_i_3_n_0),
        .O(g6371));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    g689_i_2
       (.I0(g714),
        .I1(g698),
        .I2(g673),
        .I3(g645),
        .I4(g689_i_4_n_0),
        .O(g689_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    g689_i_3
       (.I0(g689_i_5_n_0),
        .I1(g689_i_6_n_0),
        .I2(g690),
        .I3(g706),
        .I4(g677),
        .I5(g652),
        .O(g689_i_3_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_4
       (.I0(g694),
        .I1(g710),
        .I2(g647),
        .I3(g681),
        .O(g689_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    g689_i_5
       (.I0(g635),
        .I1(g669),
        .I2(g661),
        .I3(g633),
        .I4(g730),
        .I5(g723),
        .O(g689_i_5_n_0));
  LUT4 #(
    .INIT(16'hF888)) 
    g689_i_6
       (.I0(g722),
        .I1(g734),
        .I2(g634),
        .I3(g665),
        .O(g689_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g689_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6371),
        .Q(g689));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g68_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g68));
  LUT1 #(
    .INIT(2'h1)) 
    g6_i_1
       (.I0(g9310_INST_0_i_1_n_0),
        .O(g9374));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g6_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9374),
        .Q(g6));
  LUT2 #(
    .INIT(4'hB)) 
    g7048_INST_0
       (.I0(g855),
        .I1(g944),
        .O(g7048));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g706_i_1
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g706_i_2_n_0),
        .O(g706_i_1_n_0));
  LUT4 #(
    .INIT(16'hFDFF)) 
    g706_i_2
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g706_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g706_reg
       (.C(blif_clk_net),
        .CE(g706_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g706));
  LUT2 #(
    .INIT(4'h1)) 
    g7103_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7103));
  LUT4 #(
    .INIT(16'h0001)) 
    g7103_INST_0_i_1
       (.I0(g962),
        .I1(g963),
        .I2(g970),
        .I3(g7103_INST_0_i_2_n_0),
        .O(g7103_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g7103_INST_0_i_2
       (.I0(g972),
        .I1(g971),
        .I2(g966),
        .I3(g969),
        .O(g7103_INST_0_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g710_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g710));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g714_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g714));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g718_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g718));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g71_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g71));
  LUT3 #(
    .INIT(8'h6A)) 
    g727_i_1
       (.I0(g727),
        .I1(g1549),
        .I2(g1549_i_2_n_0),
        .O(g8228));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g727_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8228),
        .Q(g727));
  LUT2 #(
    .INIT(4'hB)) 
    g7283_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g7),
        .O(g7283));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    g7283_INST_0_i_1
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g58),
        .O(g7283_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g7283_INST_0_i_2
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g7283_INST_0_i_2_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g7284_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g6),
        .O(g7284));
  LUT2 #(
    .INIT(4'hB)) 
    g7285_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g5),
        .O(g7285));
  LUT2 #(
    .INIT(4'hB)) 
    g7286_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g4),
        .O(g7286));
  LUT2 #(
    .INIT(4'hB)) 
    g7287_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g2),
        .O(g7287));
  LUT2 #(
    .INIT(4'hB)) 
    g7288_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g3),
        .O(g7288));
  LUT2 #(
    .INIT(4'hB)) 
    g7289_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g48),
        .O(g7289));
  LUT2 #(
    .INIT(4'hB)) 
    g7290_INST_0
       (.I0(g7283_INST_0_i_1_n_0),
        .I1(g8),
        .O(g7290));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7291_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g48),
        .O(g7291));
  LUT5 #(
    .INIT(32'h80000000)) 
    g7291_INST_0_i_1
       (.I0(g58),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g7291_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7292_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g3),
        .O(g7292));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7293_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g2),
        .O(g7293));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    g7295_INST_0
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g4),
        .O(g7295));
  LUT2 #(
    .INIT(4'h2)) 
    g7298_INST_0
       (.I0(g1),
        .I1(g7103_INST_0_i_1_n_0),
        .O(g7298));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g730_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g730));
  LUT5 #(
    .INIT(32'h00000200)) 
    g734_i_1
       (.I0(g7291_INST_0_i_1_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .O(g734_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g734_reg
       (.C(blif_clk_net),
        .CE(g734_i_1_n_0),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g734));
  LUT6 #(
    .INIT(64'hACACACACACAFACAC)) 
    g741_i_1
       (.I0(g3),
        .I1(g741),
        .I2(g741_i_2_n_0),
        .I3(g741_i_3_n_0),
        .I4(g7480),
        .I5(g44),
        .O(g9386));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    g741_i_2
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .I4(g58),
        .I5(g746_i_2_n_0),
        .O(g741_i_2_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    g741_i_3
       (.I0(g45),
        .I1(g42),
        .I2(g41),
        .O(g741_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g741_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9386),
        .Q(g741));
  LUT6 #(
    .INIT(64'hFB08FBFBFB08FB08)) 
    g746_i_1
       (.I0(g48),
        .I1(g7291_INST_0_i_1_n_0),
        .I2(g746_i_2_n_0),
        .I3(g746),
        .I4(g741_i_3_n_0),
        .I5(g55),
        .O(g8956));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g746_i_2
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .O(g746_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g746_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8956),
        .Q(g746));
  LUT3 #(
    .INIT(8'hAB)) 
    g7474_INST_0
       (.I0(g45),
        .I1(g62),
        .I2(g65),
        .O(g7474));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g74_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g74));
  LUT4 #(
    .INIT(16'h8AAA)) 
    g7514_INST_0
       (.I0(g1034),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g7514));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g758_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g759_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g759));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g760_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g760));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g761_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g761));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g762_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g762));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g763_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g763));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g764_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g764));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g765_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g765));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g766_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g766));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g767_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8),
        .Q(g767));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g768_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g768));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g769_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g769));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g770_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g770));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g771_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g771));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g772_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g772));
  LUT2 #(
    .INIT(4'hE)) 
    g7731_INST_0
       (.I0(g16),
        .I1(g1189),
        .O(g7731));
  LUT1 #(
    .INIT(2'h1)) 
    g7732_INST_0
       (.I0(g1486),
        .O(g6223));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g773_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g3),
        .Q(g773));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g774_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g48),
        .Q(g774));
  LUT3 #(
    .INIT(8'h28)) 
    g775_i_1
       (.I0(g781),
        .I1(g775_i_2_n_0),
        .I2(g775),
        .O(g7759));
  LUT5 #(
    .INIT(32'h80000000)) 
    g775_i_2
       (.I0(g812),
        .I1(g806),
        .I2(g799),
        .I3(g803),
        .I4(g809),
        .O(g775_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g775_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7759),
        .Q(g775));
  LUT2 #(
    .INIT(4'h6)) 
    g778_i_1
       (.I0(g778),
        .I1(g778_i_2_n_0),
        .O(g7296));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g778_i_2
       (.I0(g809),
        .I1(g803),
        .I2(g799),
        .I3(g806),
        .I4(g812),
        .I5(g775),
        .O(g778_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g778_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7296),
        .Q(g778));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g77_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g77));
  LUT3 #(
    .INIT(8'h6A)) 
    g782_i_1
       (.I0(g782),
        .I1(g792),
        .I2(g795),
        .O(g5734));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g782_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5734),
        .Q(g782));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    g786_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g815),
        .I3(g819),
        .I4(g822),
        .I5(g828),
        .O(g786_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g786_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g786_i_1_n_0),
        .Q(g786));
  LUT2 #(
    .INIT(4'h6)) 
    g789_i_1
       (.I0(g789),
        .I1(g5287),
        .O(g7297));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    g789_i_2
       (.I0(g828),
        .I1(g822),
        .I2(g819),
        .I3(g815),
        .I4(g825),
        .I5(g786),
        .O(g5287));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g789_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7297),
        .Q(g789));
  LUT2 #(
    .INIT(4'h6)) 
    g792_i_1
       (.I0(g792),
        .I1(g795),
        .O(g792_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g792_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g792_i_1_n_0),
        .Q(g792));
  LUT1 #(
    .INIT(2'h1)) 
    g795_i_1
       (.I0(g795),
        .O(g1683));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g795_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1683),
        .Q(g795));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .O(g7756));
  LUT2 #(
    .INIT(4'h2)) 
    g799_i_2
       (.I0(g781),
        .I1(g778_i_2_n_0),
        .O(g799_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g799_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7756),
        .Q(g799));
  LUT1 #(
    .INIT(2'h1)) 
    g7_i_1
       (.I0(g9312_INST_0_i_1_n_0),
        .O(g9375));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g7_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9375),
        .Q(g7));
  LUT3 #(
    .INIT(8'h28)) 
    g803_i_1
       (.I0(g799_i_2_n_0),
        .I1(g799),
        .I2(g803),
        .O(g7757));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g803_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7757),
        .Q(g803));
  LUT4 #(
    .INIT(16'h78FF)) 
    g806_i_1
       (.I0(g803),
        .I1(g799),
        .I2(g806),
        .I3(g799_i_2_n_0),
        .O(g7510));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g806_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7510),
        .Q(g806));
  LUT5 #(
    .INIT(32'h7F80FFFF)) 
    g809_i_1
       (.I0(g806),
        .I1(g799),
        .I2(g803),
        .I3(g809),
        .I4(g799_i_2_n_0),
        .O(g7511));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g809_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7511),
        .Q(g809));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g80_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g80));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    g812_i_1
       (.I0(g799_i_2_n_0),
        .I1(g809),
        .I2(g803),
        .I3(g799),
        .I4(g806),
        .I5(g812),
        .O(g7758));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g812_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7758),
        .Q(g812));
  LUT1 #(
    .INIT(2'h1)) 
    g815_i_1
       (.I0(g815),
        .O(g815_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g815_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g815_i_1_n_0),
        .Q(g815));
  LUT2 #(
    .INIT(4'h6)) 
    g819_i_1
       (.I0(g815),
        .I1(g819),
        .O(g819_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g819_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g819_i_1_n_0),
        .Q(g819));
  LUT1 #(
    .INIT(2'h1)) 
    g8219_INST_0
       (.I0(g1432),
        .O(g6675));
  LUT6 #(
    .INIT(64'h80FFFF00FF00FF00)) 
    g822_i_1
       (.I0(g786),
        .I1(g825),
        .I2(g828),
        .I3(g822),
        .I4(g815),
        .I5(g819),
        .O(g822_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g822_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g822_i_1_n_0),
        .Q(g822));
  LUT6 #(
    .INIT(64'h8FF0F0F0F0F0F0F0)) 
    g825_i_1
       (.I0(g786),
        .I1(g828),
        .I2(g825),
        .I3(g822),
        .I4(g819),
        .I5(g815),
        .O(g825_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g825_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g825_i_1_n_0),
        .Q(g825));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    g828_i_1
       (.I0(g825),
        .I1(g815),
        .I2(g819),
        .I3(g822),
        .I4(g828),
        .O(g828_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g828_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g828_i_1_n_0),
        .Q(g828));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g831_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g831));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g834_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g834));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g837_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g837));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g83_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6),
        .Q(g83));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g840_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g840));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g843_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g843));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g846_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g846));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g849_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g849));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g852_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g883),
        .Q(g852));
  LUT3 #(
    .INIT(8'hB8)) 
    g855_i_1
       (.I0(g48),
        .I1(g859_i_2_n_0),
        .I2(g855),
        .O(g8220));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g855_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8220),
        .Q(g855));
  LUT3 #(
    .INIT(8'hB8)) 
    g859_i_1
       (.I0(g3),
        .I1(g859_i_2_n_0),
        .I2(g859),
        .O(g8221));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    g859_i_2
       (.I0(g58),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g859_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g859_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8221),
        .Q(g859));
  LUT4 #(
    .INIT(16'hBBB8)) 
    g863_i_1
       (.I0(g2),
        .I1(g859_i_2_n_0),
        .I2(g866),
        .I3(g863),
        .O(g8222));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g863_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8222),
        .Q(g863));
  LUT2 #(
    .INIT(4'h7)) 
    g8663_INST_0
       (.I0(g1412),
        .I1(g1405),
        .O(g8663));
  LUT2 #(
    .INIT(4'h2)) 
    g866_i_1
       (.I0(g874),
        .I1(g878),
        .O(g5163));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g866_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5163),
        .Q(g866));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g86_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7),
        .Q(g86));
  LUT3 #(
    .INIT(8'h6A)) 
    g871_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g5167));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g871_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5167),
        .Q(g871));
  LUT3 #(
    .INIT(8'h80)) 
    g874_i_1
       (.I0(g871),
        .I1(g929),
        .I2(g933),
        .O(g4654));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g874_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4654),
        .Q(g874));
  LUT4 #(
    .INIT(16'h0080)) 
    g875_i_1
       (.I0(g878),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g5165));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g875_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5165),
        .Q(g875));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g878_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g890),
        .Q(g878));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g883_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g921),
        .Q(g883));
  LUT3 #(
    .INIT(8'h4F)) 
    g8872_INST_0
       (.I0(g1030),
        .I1(g8872_INST_0_i_1_n_0),
        .I2(g1),
        .O(g8872));
  LUT4 #(
    .INIT(16'h4555)) 
    g8872_INST_0_i_1
       (.I0(g7566),
        .I1(g979),
        .I2(g43),
        .I3(g984),
        .O(g8872_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0CFC0CCCCCFFCCCE)) 
    g887_i_1
       (.I0(g887_i_2_n_0),
        .I1(g887),
        .I2(g889),
        .I3(g888),
        .I4(g926),
        .I5(g4654),
        .O(g7099));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    g887_i_2
       (.I0(g866),
        .I1(g887_i_3_n_0),
        .I2(g896),
        .I3(g906),
        .I4(g901),
        .I5(g883),
        .O(g887_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g887_i_3
       (.I0(g921),
        .I1(g911),
        .I2(g916),
        .I3(g891),
        .O(g887_i_3_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g887_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7099),
        .Q(g887));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAEAEAEA)) 
    g888_i_1
       (.I0(g888_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g875),
        .O(g7100));
  LUT5 #(
    .INIT(32'h000A0030)) 
    g888_i_2
       (.I0(g866),
        .I1(g878),
        .I2(g887),
        .I3(g888),
        .I4(g889),
        .O(g888_i_2_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g888_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7100),
        .Q(g888));
  LUT6 #(
    .INIT(64'hBAAAFAAAAAAAEAAA)) 
    g889_i_1
       (.I0(g889_i_2_n_0),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .I4(g4654),
        .I5(g874),
        .O(g7101));
  LUT6 #(
    .INIT(64'h5555555445444544)) 
    g889_i_2
       (.I0(g926),
        .I1(g889_i_3_n_0),
        .I2(g866),
        .I3(g889_i_4_n_0),
        .I4(g889_i_5_n_0),
        .I5(g889_i_6_n_0),
        .O(g889_i_2_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    g889_i_3
       (.I0(g888),
        .I1(g889),
        .I2(g887),
        .O(g889_i_3_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    g889_i_4
       (.I0(g875),
        .I1(g888),
        .I2(g887),
        .I3(g889),
        .O(g889_i_4_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    g889_i_5
       (.I0(g883),
        .I1(g901),
        .I2(g906),
        .I3(g896),
        .I4(g887_i_3_n_0),
        .O(g889_i_5_n_0));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    g889_i_6
       (.I0(g933),
        .I1(g929),
        .I2(g871),
        .I3(g888),
        .I4(g889),
        .I5(g887),
        .O(g889_i_6_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g889_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7101),
        .Q(g889));
  LUT3 #(
    .INIT(8'hB8)) 
    g890_i_1
       (.I0(g12),
        .I1(g859),
        .I2(g11),
        .O(g7102));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g890_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7102),
        .Q(g890));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g891_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g926),
        .Q(g891));
  LUT6 #(
    .INIT(64'hAAAAAAAA2000AAAA)) 
    g8958_INST_0
       (.I0(g8872),
        .I1(g1029),
        .I2(g1033),
        .I3(g43),
        .I4(g1),
        .I5(g10),
        .O(g8958));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g896_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g891),
        .Q(g896));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g89_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g92),
        .Q(g89));
  (* KEEP = "yes" *) 
  FDCE #(
    .INIT(1'b0)) 
    g8_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9376),
        .Q(g8));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g901_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g896),
        .Q(g901));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g906_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g901),
        .Q(g906));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g911_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g906),
        .Q(g911));
  LUT3 #(
    .INIT(8'hF7)) 
    g9132_INST_0
       (.I0(g43),
        .I1(g1033),
        .I2(g1029),
        .O(g9132));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g916_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g911),
        .Q(g916));
  LUT3 #(
    .INIT(8'hB8)) 
    g9204_INST_0
       (.I0(g30),
        .I1(g32),
        .I2(g31),
        .O(g9204));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g921_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g916),
        .Q(g921));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g926_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g878),
        .Q(g926));
  LUT2 #(
    .INIT(4'h7)) 
    g9280_INST_0
       (.I0(g62),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9280));
  LUT6 #(
    .INIT(64'hFF10FF10FFFFFF10)) 
    g9280_INST_0_i_1
       (.I0(g9280_INST_0_i_2_n_0),
        .I1(g9280_INST_0_i_3_n_0),
        .I2(g9280_INST_0_i_4_n_0),
        .I3(g9280_INST_0_i_5_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9280_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_10
       (.I0(g632),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    g9280_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9280_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_12
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g110),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_33_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g228),
        .O(g9280_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g553),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g365),
        .O(g9280_INST_0_i_13_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_14
       (.I0(g608),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_25_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9280_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    g9280_INST_0_i_15
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9280_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9280_INST_0_i_16
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g284),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g185),
        .O(g9280_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_17
       (.I0(g746_i_2_n_0),
        .I1(g446),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g309),
        .O(g9280_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    g9280_INST_0_i_18
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9280_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_19
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9280_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9280_INST_0_i_2
       (.I0(g9280_INST_0_i_8_n_0),
        .I1(g9280_INST_0_i_9_n_0),
        .I2(g9280_INST_0_i_10_n_0),
        .I3(g9280_INST_0_i_11_n_0),
        .I4(g613),
        .I5(g9280_INST_0_i_12_n_0),
        .O(g9280_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_20
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g855),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g852),
        .O(g9280_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0C0CFF0C0C0CAEAE)) 
    g9280_INST_0_i_21
       (.I0(g758),
        .I1(g774),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g766),
        .I4(g9305_INST_0_i_27_n_0),
        .I5(g68),
        .O(g9280_INST_0_i_21_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    g9280_INST_0_i_22
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .O(g9280_INST_0_i_22_n_0));
  LUT4 #(
    .INIT(16'hF8D9)) 
    g9280_INST_0_i_23
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9280_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    g9280_INST_0_i_24
       (.I0(g52),
        .I1(g80),
        .I2(g86),
        .I3(g83),
        .O(g9280_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_25
       (.I0(g746),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g746_i_2_n_0),
        .O(g9280_INST_0_i_25_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_26
       (.I0(g527),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9280_INST_0_i_26_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_27
       (.I0(g471),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9280_INST_0_i_27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9280_INST_0_i_28
       (.I0(g694),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9280_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g685),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g648),
        .O(g9280_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    g9280_INST_0_i_3
       (.I0(g9280_INST_0_i_13_n_0),
        .I1(g9280_INST_0_i_14_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g621),
        .I4(g9280_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_17_n_0),
        .O(g9280_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9280_INST_0_i_30
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g49),
        .I2(g9280_INST_0_i_32_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g710),
        .O(g9280_INST_0_i_30_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_31
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .O(g9280_INST_0_i_31_n_0));
  LUT4 #(
    .INIT(16'hFFFB)) 
    g9280_INST_0_i_32
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    g9280_INST_0_i_33
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9280_INST_0_i_33_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9280_INST_0_i_34
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .O(g9280_INST_0_i_34_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_35
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9280_INST_0_i_35_n_0));
  LUT4 #(
    .INIT(16'hFBFF)) 
    g9280_INST_0_i_36
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9280_INST_0_i_36_n_0));
  LUT4 #(
    .INIT(16'hB0BB)) 
    g9280_INST_0_i_4
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g142),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g168),
        .O(g9280_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h4500450000004500)) 
    g9280_INST_0_i_5
       (.I0(g9280_INST_0_i_20_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g48),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_21_n_0),
        .I5(g498_i_2_n_0),
        .O(g9280_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000111100001FFF)) 
    g9280_INST_0_i_6
       (.I0(g9280_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_23_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g9280_INST_0_i_24_n_0),
        .O(g9280_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9280_INST_0_i_7
       (.I0(g9280_INST_0_i_25_n_0),
        .I1(g9280_INST_0_i_26_n_0),
        .I2(g9280_INST_0_i_27_n_0),
        .I3(g9280_INST_0_i_28_n_0),
        .I4(g9280_INST_0_i_29_n_0),
        .I5(g9280_INST_0_i_30_n_0),
        .O(g9280_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFCF8FCFFFCF8FCF0)) 
    g9280_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g624),
        .O(g9280_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9280_INST_0_i_9
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g600),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g390),
        .O(g9280_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9297_INST_0
       (.I0(g9360),
        .I1(g62),
        .O(g9297));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    g9297_INST_0_i_1
       (.I0(g9297_INST_0_i_2_n_0),
        .I1(g9297_INST_0_i_3_n_0),
        .I2(g9297_INST_0_i_4_n_0),
        .I3(g9297_INST_0_i_5_n_0),
        .I4(g9297_INST_0_i_6_n_0),
        .I5(g9297_INST_0_i_7_n_0),
        .O(g9360));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_10
       (.I0(g746_i_2_n_0),
        .I1(g443),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_29_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g362),
        .O(g9297_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9297_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9297_INST_0_i_12
       (.I0(g631),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9297_INST_0_i_13
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g182),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g162),
        .O(g9297_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_14
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g281),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_36_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g306),
        .O(g9297_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9297_INST_0_i_15
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g225),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g607),
        .O(g9297_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9297_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g68),
        .I3(g77),
        .I4(g74),
        .I5(g71),
        .O(g9297_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9297_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_18
       (.I0(g105),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9297_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_19
       (.I0(g9299_INST_0_i_29_n_0),
        .I1(g859),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g849),
        .O(g9297_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    g9297_INST_0_i_2
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g599),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9297_INST_0_i_9_n_0),
        .I4(g68),
        .I5(g612),
        .O(g9297_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFB0FFFFFFBB)) 
    g9297_INST_0_i_20
       (.I0(g706_i_2_n_0),
        .I1(g765),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g773),
        .O(g9297_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_21
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g714),
        .I2(g9305_INST_0_i_7_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g698),
        .O(g9297_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_22
       (.I0(g746_i_2_n_0),
        .I1(g741),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g647),
        .O(g9297_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9297_INST_0_i_23
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g757),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g681),
        .O(g9297_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000000E00000002)) 
    g9297_INST_0_i_24
       (.I0(g468),
        .I1(g68),
        .I2(g9280_INST_0_i_22_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g524),
        .O(g9297_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    g9297_INST_0_i_3
       (.I0(g9297_INST_0_i_10_n_0),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g550),
        .I3(g9297_INST_0_i_12_n_0),
        .I4(g9297_INST_0_i_13_n_0),
        .I5(g9297_INST_0_i_14_n_0),
        .O(g9297_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9297_INST_0_i_4
       (.I0(g9297_INST_0_i_15_n_0),
        .I1(g623),
        .I2(g9297_INST_0_i_16_n_0),
        .I3(g620),
        .I4(g9280_INST_0_i_15_n_0),
        .O(g9297_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2F2FFF2)) 
    g9297_INST_0_i_5
       (.I0(g138),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g387),
        .I4(g9297_INST_0_i_17_n_0),
        .I5(g9297_INST_0_i_18_n_0),
        .O(g9297_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h45000000)) 
    g9297_INST_0_i_6
       (.I0(g9297_INST_0_i_19_n_0),
        .I1(g9299_INST_0_i_12_n_0),
        .I2(g3),
        .I3(g9297_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_4_n_0),
        .O(g9297_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9297_INST_0_i_7
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9297_INST_0_i_21_n_0),
        .I2(g9297_INST_0_i_22_n_0),
        .I3(g9297_INST_0_i_23_n_0),
        .I4(g9297_INST_0_i_24_n_0),
        .O(g9297_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    g9297_INST_0_i_8
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9297_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    g9297_INST_0_i_9
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .O(g9297_INST_0_i_9_n_0));
  LUT6 #(
    .INIT(64'h00005155FFFFFFFF)) 
    g9299_INST_0
       (.I0(g9299_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_3_n_0),
        .I3(g9299_INST_0_i_4_n_0),
        .I4(g9299_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9299));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    g9299_INST_0_i_1
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9299_INST_0_i_6_n_0),
        .I2(g9299_INST_0_i_7_n_0),
        .I3(g9299_INST_0_i_8_n_0),
        .I4(g9299_INST_0_i_9_n_0),
        .I5(g9299_INST_0_i_10_n_0),
        .O(g9299_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02023302)) 
    g9299_INST_0_i_10
       (.I0(g134),
        .I1(g573_i_2_n_0),
        .I2(g706_i_2_n_0),
        .I3(g351),
        .I4(g9299_INST_0_i_29_n_0),
        .I5(g9299_INST_0_i_30_n_0),
        .O(g9299_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    g9299_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g68),
        .O(g9299_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_12
       (.I0(g68),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    g9299_INST_0_i_13
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    g9299_INST_0_i_14
       (.I0(g68),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    g9299_INST_0_i_15
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_15_n_0));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    g9299_INST_0_i_16
       (.I0(g41),
        .I1(g42),
        .I2(g45),
        .I3(g44),
        .I4(g55),
        .O(g9299_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9299_INST_0_i_17
       (.I0(g52),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .O(g9299_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9299_INST_0_i_18
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g702),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g677),
        .O(g9299_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    g9299_INST_0_i_19
       (.I0(g513),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9299_INST_0_i_2
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9299_INST_0_i_12_n_0),
        .I4(g846),
        .I5(g9299_INST_0_i_13_n_0),
        .O(g9299_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_20
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9299_INST_0_i_21
       (.I0(g718),
        .I1(g9299_INST_0_i_31_n_0),
        .I2(g465),
        .I3(g9305_INST_0_i_20_n_0),
        .I4(g9299_INST_0_i_32_n_0),
        .I5(g756),
        .O(g9299_INST_0_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9299_INST_0_i_22
       (.I0(g222),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9299_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_23
       (.I0(g9305_INST_0_i_28_n_0),
        .I1(g598),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g181),
        .O(g9299_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9299_INST_0_i_24
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'h444F4444)) 
    g9299_INST_0_i_25
       (.I0(g4_i_3_n_0),
        .I1(g100),
        .I2(g746_i_2_n_0),
        .I3(g573_i_2_n_0),
        .I4(g432),
        .O(g9299_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g9299_INST_0_i_26
       (.I0(g630),
        .I1(g498_i_2_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9299_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9299_INST_0_i_27
       (.I0(g611),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9299_INST_0_i_27_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    g9299_INST_0_i_28
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9299_INST_0_i_28_n_0));
  LUT4 #(
    .INIT(16'hDFFF)) 
    g9299_INST_0_i_29
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g68),
        .O(g9299_INST_0_i_29_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9299_INST_0_i_3
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g764),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g772),
        .O(g9299_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9299_INST_0_i_30
       (.I0(g9305_INST_0_i_25_n_0),
        .I1(g606),
        .I2(g9280_INST_0_i_34_n_0),
        .I3(g573_i_2_n_0),
        .I4(g547),
        .O(g9299_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_31
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9299_INST_0_i_32
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9299_INST_0_i_32_n_0));
  LUT5 #(
    .INIT(32'h0000003E)) 
    g9299_INST_0_i_4
       (.I0(g71),
        .I1(g77),
        .I2(g74),
        .I3(g9299_INST_0_i_16_n_0),
        .I4(g9299_INST_0_i_17_n_0),
        .O(g9299_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    g9299_INST_0_i_5
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_18_n_0),
        .I2(g9299_INST_0_i_19_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .I5(g9299_INST_0_i_21_n_0),
        .O(g9299_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    g9299_INST_0_i_6
       (.I0(g9299_INST_0_i_17_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g9305_INST_0_i_6_n_0),
        .O(g9299_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h1011000010111011)) 
    g9299_INST_0_i_7
       (.I0(g9299_INST_0_i_22_n_0),
        .I1(g9299_INST_0_i_23_n_0),
        .I2(g9299_INST_0_i_24_n_0),
        .I3(g270),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g619),
        .O(g9299_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFAAAEAAAEAAAE)) 
    g9299_INST_0_i_8
       (.I0(g9299_INST_0_i_25_n_0),
        .I1(g622),
        .I2(g498_i_2_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g384),
        .I5(g573_i_1_n_0),
        .O(g9299_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    g9299_INST_0_i_9
       (.I0(g9299_INST_0_i_26_n_0),
        .I1(g9299_INST_0_i_27_n_0),
        .I2(g158),
        .I3(g9299_INST_0_i_28_n_0),
        .I4(g303),
        .I5(g9305_INST_0_i_8_n_0),
        .O(g9299_INST_0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    g929_i_1
       (.I0(g929),
        .O(g1681));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g929_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1681),
        .Q(g929));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g92_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5),
        .Q(g92));
  LUT6 #(
    .INIT(64'h0000FE00FFFFFFFF)) 
    g9305_INST_0
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9305_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_3_n_0),
        .I3(g9305_INST_0_i_4_n_0),
        .I4(g9305_INST_0_i_5_n_0),
        .I5(g62),
        .O(g9305));
  LUT5 #(
    .INIT(32'hEEECECEC)) 
    g9305_INST_0_i_1
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .O(g9305_INST_0_i_1_n_0));
  LUT5 #(
    .INIT(32'h004F0044)) 
    g9305_INST_0_i_10
       (.I0(g706_i_2_n_0),
        .I1(g130),
        .I2(g9299_INST_0_i_29_n_0),
        .I3(g573_i_2_n_0),
        .I4(g348),
        .O(g9305_INST_0_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    g9305_INST_0_i_11
       (.I0(g219),
        .I1(g9305_INST_0_i_23_n_0),
        .O(g9305_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF004400F4)) 
    g9305_INST_0_i_12
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g154),
        .I2(g180),
        .I3(g573_i_2_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g9305_INST_0_i_24_n_0),
        .O(g9305_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8)) 
    g9305_INST_0_i_13
       (.I0(g381),
        .I1(g573_i_1_n_0),
        .I2(g605),
        .I3(g573_i_2_n_0),
        .I4(g9305_INST_0_i_25_n_0),
        .I5(g9305_INST_0_i_26_n_0),
        .O(g9305_INST_0_i_13_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9305_INST_0_i_14
       (.I0(g95),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_27_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_15
       (.I0(g573_i_2_n_0),
        .I1(g68),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .O(g9305_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h101010FF10101010)) 
    g9305_INST_0_i_16
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g629),
        .I3(g9305_INST_0_i_28_n_0),
        .I4(g573_i_2_n_0),
        .I5(g597),
        .O(g9305_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9305_INST_0_i_17
       (.I0(g9299_INST_0_i_20_n_0),
        .I1(g645),
        .I2(g753),
        .I3(g9299_INST_0_i_32_n_0),
        .I4(g673),
        .I5(g9305_INST_0_i_29_n_0),
        .O(g9305_INST_0_i_17_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_18
       (.I0(g9305_INST_0_i_30_n_0),
        .I1(g510),
        .I2(g9305_INST_0_i_31_n_0),
        .I3(g722),
        .O(g9305_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    g9305_INST_0_i_19
       (.I0(g734),
        .I1(g9305_INST_0_i_32_n_0),
        .I2(g68),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF5D)) 
    g9305_INST_0_i_2
       (.I0(g9299_INST_0_i_6_n_0),
        .I1(g300),
        .I2(g9305_INST_0_i_8_n_0),
        .I3(g9305_INST_0_i_9_n_0),
        .I4(g9305_INST_0_i_10_n_0),
        .I5(g9305_INST_0_i_11_n_0),
        .O(g9305_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    g9305_INST_0_i_20
       (.I0(g71),
        .I1(g74),
        .I2(g77),
        .I3(g68),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_20_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9305_INST_0_i_21
       (.I0(g9299_INST_0_i_14_n_0),
        .I1(g763),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g771),
        .O(g9305_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    g9305_INST_0_i_22
       (.I0(g68),
        .I1(g55),
        .I2(g44),
        .I3(g45),
        .I4(g42),
        .I5(g41),
        .O(g9305_INST_0_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    g9305_INST_0_i_23
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_23_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9305_INST_0_i_24
       (.I0(g267),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9280_INST_0_i_35_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_24_n_0));
  LUT4 #(
    .INIT(16'hF7FF)) 
    g9305_INST_0_i_25
       (.I0(g77),
        .I1(g74),
        .I2(g71),
        .I3(g68),
        .O(g9305_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000C0800000008)) 
    g9305_INST_0_i_26
       (.I0(g429),
        .I1(g68),
        .I2(g9305_INST_0_i_33_n_0),
        .I3(g71),
        .I4(g573_i_2_n_0),
        .I5(g573),
        .O(g9305_INST_0_i_26_n_0));
  LUT3 #(
    .INIT(8'hEF)) 
    g9305_INST_0_i_27
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9305_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'hFFBF)) 
    g9305_INST_0_i_28
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_29
       (.I0(g706_i_2_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    g9305_INST_0_i_3
       (.I0(g9305_INST_0_i_12_n_0),
        .I1(g9305_INST_0_i_13_n_0),
        .I2(g9305_INST_0_i_14_n_0),
        .I3(g618),
        .I4(g9305_INST_0_i_15_n_0),
        .I5(g9305_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    g9305_INST_0_i_30
       (.I0(g68),
        .I1(g71),
        .I2(g74),
        .I3(g77),
        .I4(g9299_INST_0_i_17_n_0),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    g9305_INST_0_i_31
       (.I0(g9305_INST_0_i_7_n_0),
        .I1(g52),
        .I2(g80),
        .I3(g86),
        .I4(g83),
        .I5(g9299_INST_0_i_16_n_0),
        .O(g9305_INST_0_i_31_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    g9305_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g83),
        .I2(g86),
        .I3(g80),
        .I4(g52),
        .O(g9305_INST_0_i_32_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9305_INST_0_i_33
       (.I0(g74),
        .I1(g77),
        .O(g9305_INST_0_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFFFEFFFFFFFF)) 
    g9305_INST_0_i_4
       (.I0(g9305_INST_0_i_17_n_0),
        .I1(g9305_INST_0_i_18_n_0),
        .I2(g9305_INST_0_i_19_n_0),
        .I3(g462),
        .I4(g9305_INST_0_i_20_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9305_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9305_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9305_INST_0_i_21_n_0),
        .I2(g9299_INST_0_i_12_n_0),
        .I3(g4),
        .I4(g9299_INST_0_i_13_n_0),
        .I5(g843),
        .O(g9305_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_6
       (.I0(g80),
        .I1(g52),
        .I2(g83),
        .I3(g86),
        .O(g9305_INST_0_i_6_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    g9305_INST_0_i_7
       (.I0(g68),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .O(g9305_INST_0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    g9305_INST_0_i_8
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .I3(g68),
        .I4(g573_i_2_n_0),
        .O(g9305_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    g9305_INST_0_i_9
       (.I0(g610),
        .I1(g9305_INST_0_i_22_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g71),
        .I4(g77),
        .I5(g74),
        .O(g9305_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9308_INST_0
       (.I0(g62),
        .I1(g9308_INST_0_i_1_n_0),
        .O(g9308));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    g9308_INST_0_i_1
       (.I0(g9308_INST_0_i_2_n_0),
        .I1(g9308_INST_0_i_3_n_0),
        .I2(g9305_INST_0_i_1_n_0),
        .I3(g9308_INST_0_i_4_n_0),
        .I4(g9280_INST_0_i_6_n_0),
        .I5(g9308_INST_0_i_5_n_0),
        .O(g9308_INST_0_i_1_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_10
       (.I0(g628),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'h00000200)) 
    g9308_INST_0_i_11
       (.I0(g617),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000002300000020)) 
    g9308_INST_0_i_12
       (.I0(g345),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g9308_INST_0_i_24_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g297),
        .O(g9308_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_13
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g591),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g426),
        .O(g9308_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9308_INST_0_i_14
       (.I0(g706_i_2_n_0),
        .I1(g126),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9305_INST_0_i_7_n_0),
        .I5(g174),
        .O(g9308_INST_0_i_14_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_15
       (.I0(g179),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_16
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g840),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g5),
        .O(g9308_INST_0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_17
       (.I0(g507),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .O(g9308_INST_0_i_17_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_18
       (.I0(g730),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g68),
        .I4(g9305_INST_0_i_27_n_0),
        .O(g9308_INST_0_i_18_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_19
       (.I0(g459),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_28_n_0),
        .O(g9308_INST_0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_2
       (.I0(g9308_INST_0_i_6_n_0),
        .I1(g9308_INST_0_i_7_n_0),
        .I2(g9308_INST_0_i_8_n_0),
        .I3(g9308_INST_0_i_9_n_0),
        .I4(g9308_INST_0_i_10_n_0),
        .I5(g9308_INST_0_i_11_n_0),
        .O(g9308_INST_0_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_20
       (.I0(g723),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9308_INST_0_i_20_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9308_INST_0_i_21
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g752),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g669),
        .O(g9308_INST_0_i_21_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_22
       (.I0(g635),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9280_INST_0_i_24_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9308_INST_0_i_22_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    g9308_INST_0_i_23
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_23_n_0));
  LUT3 #(
    .INIT(8'hDF)) 
    g9308_INST_0_i_24
       (.I0(g74),
        .I1(g77),
        .I2(g71),
        .O(g9308_INST_0_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    g9308_INST_0_i_3
       (.I0(g9308_INST_0_i_12_n_0),
        .I1(g9308_INST_0_i_13_n_0),
        .I2(g9308_INST_0_i_14_n_0),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g264),
        .I5(g9308_INST_0_i_15_n_0),
        .O(g9308_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9308_INST_0_i_4
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9308_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g762),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g770),
        .O(g9308_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g9308_INST_0_i_5
       (.I0(g9308_INST_0_i_17_n_0),
        .I1(g9308_INST_0_i_18_n_0),
        .I2(g9308_INST_0_i_19_n_0),
        .I3(g9308_INST_0_i_20_n_0),
        .I4(g9308_INST_0_i_21_n_0),
        .I5(g9308_INST_0_i_22_n_0),
        .O(g9308_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_6
       (.I0(g9280_INST_0_i_33_n_0),
        .I1(g216),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g378),
        .O(g9308_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9308_INST_0_i_7
       (.I0(g9280_INST_0_i_32_n_0),
        .I1(g89),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g604),
        .O(g9308_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9308_INST_0_i_8
       (.I0(g596),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g9305_INST_0_i_28_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'h00000002)) 
    g9308_INST_0_i_9
       (.I0(g609),
        .I1(g68),
        .I2(g9308_INST_0_i_23_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .O(g9308_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9310_INST_0
       (.I0(g62),
        .I1(g9310_INST_0_i_1_n_0),
        .O(g9310));
  LUT6 #(
    .INIT(64'h00000F00EEEEEEEE)) 
    g9310_INST_0_i_1
       (.I0(g9310_INST_0_i_2_n_0),
        .I1(g9310_INST_0_i_3_n_0),
        .I2(g9310_INST_0_i_4_n_0),
        .I3(g9310_INST_0_i_5_n_0),
        .I4(g9310_INST_0_i_6_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9310_INST_0_i_10
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g261),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g423),
        .O(g9310_INST_0_i_10_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9310_INST_0_i_11
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g706_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g122),
        .O(g9310_INST_0_i_11_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9310_INST_0_i_12
       (.I0(g627),
        .I1(g7283_INST_0_i_2_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9310_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    g9310_INST_0_i_13
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g71),
        .I2(g77),
        .I3(g74),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9310_INST_0_i_14
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9310_INST_0_i_14_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9310_INST_0_i_2
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9310_INST_0_i_7_n_0),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g769),
        .I4(g9299_INST_0_i_14_n_0),
        .I5(g761),
        .O(g9310_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9310_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g754),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g504),
        .I5(g9310_INST_0_i_8_n_0),
        .O(g9310_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9310_INST_0_i_4
       (.I0(g588),
        .I1(g9297_INST_0_i_11_n_0),
        .I2(g603),
        .I3(g9310_INST_0_i_9_n_0),
        .I4(g9310_INST_0_i_10_n_0),
        .O(g9310_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h00D000D0000000D0)) 
    g9310_INST_0_i_5
       (.I0(g616),
        .I1(g9280_INST_0_i_15_n_0),
        .I2(g9310_INST_0_i_11_n_0),
        .I3(g9310_INST_0_i_12_n_0),
        .I4(g342),
        .I5(g9310_INST_0_i_13_n_0),
        .O(g9310_INST_0_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9310_INST_0_i_6
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g184),
        .I2(g9310_INST_0_i_14_n_0),
        .I3(g150),
        .I4(g9280_INST_0_i_19_n_0),
        .O(g9310_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g837),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g6),
        .O(g9310_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9310_INST_0_i_8
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g634),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g665),
        .O(g9310_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    g9310_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g77),
        .I2(g74),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9310_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    g9312_INST_0
       (.I0(g62),
        .I1(g9312_INST_0_i_1_n_0),
        .O(g9312));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    g9312_INST_0_i_1
       (.I0(g9312_INST_0_i_2_n_0),
        .I1(g9312_INST_0_i_3_n_0),
        .I2(g9312_INST_0_i_4_n_0),
        .I3(g9312_INST_0_i_5_n_0),
        .I4(g9312_INST_0_i_6_n_0),
        .I5(g9312_INST_0_i_7_n_0),
        .O(g9312_INST_0_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9312_INST_0_i_10
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g633),
        .I2(g706_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g661),
        .O(g9312_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    g9312_INST_0_i_11
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g77),
        .I3(g74),
        .I4(g71),
        .I5(g68),
        .O(g9312_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9312_INST_0_i_12
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g258),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g420),
        .O(g9312_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_2
       (.I0(g9312_INST_0_i_8_n_0),
        .I1(g9299_INST_0_i_15_n_0),
        .I2(g768),
        .I3(g9299_INST_0_i_14_n_0),
        .I4(g760),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9312_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000008A008A8A)) 
    g9312_INST_0_i_3
       (.I0(g9280_INST_0_i_6_n_0),
        .I1(g9299_INST_0_i_32_n_0),
        .I2(g755),
        .I3(g9305_INST_0_i_30_n_0),
        .I4(g501),
        .I5(g9312_INST_0_i_10_n_0),
        .O(g9312_INST_0_i_3_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9312_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g173),
        .I2(g9280_INST_0_i_19_n_0),
        .I3(g183),
        .I4(g9310_INST_0_i_14_n_0),
        .O(g9312_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    g9312_INST_0_i_5
       (.I0(g9310_INST_0_i_13_n_0),
        .I1(g339),
        .I2(g9312_INST_0_i_11_n_0),
        .I3(g626),
        .O(g9312_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'hD0DD)) 
    g9312_INST_0_i_6
       (.I0(g118),
        .I1(g9280_INST_0_i_18_n_0),
        .I2(g9280_INST_0_i_15_n_0),
        .I3(g615),
        .O(g9312_INST_0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9312_INST_0_i_7
       (.I0(g602),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g570),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9312_INST_0_i_12_n_0),
        .O(g9312_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFF0FFFDFFFD)) 
    g9312_INST_0_i_8
       (.I0(g834),
        .I1(g9280_INST_0_i_34_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g746_i_2_n_0),
        .I5(g7),
        .O(g9312_INST_0_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFEEEEEF)) 
    g9312_INST_0_i_9
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .O(g9312_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    g9314_INST_0
       (.I0(g9376),
        .I1(g62),
        .O(g9314));
  LUT6 #(
    .INIT(64'hFB00FBFFFB00FB00)) 
    g9314_INST_0_i_1
       (.I0(g9314_INST_0_i_2_n_0),
        .I1(g9314_INST_0_i_3_n_0),
        .I2(g9314_INST_0_i_4_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9314_INST_0_i_5_n_0),
        .I5(g9314_INST_0_i_6_n_0),
        .O(g9376));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_10
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g831),
        .I2(g746_i_2_n_0),
        .I3(g9299_INST_0_i_17_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g8),
        .O(g9314_INST_0_i_10_n_0));
  LUT6 #(
    .INIT(64'h0000004F00000044)) 
    g9314_INST_0_i_11
       (.I0(g706_i_2_n_0),
        .I1(g706),
        .I2(g7283_INST_0_i_2_n_0),
        .I3(g9280_INST_0_i_24_n_0),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g690),
        .O(g9314_INST_0_i_11_n_0));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    g9314_INST_0_i_2
       (.I0(g336),
        .I1(g9310_INST_0_i_13_n_0),
        .I2(g255),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g9314_INST_0_i_7_n_0),
        .O(g9314_INST_0_i_2_n_0));
  LUT6 #(
    .INIT(64'h00000000D0D000D0)) 
    g9314_INST_0_i_3
       (.I0(g625),
        .I1(g9312_INST_0_i_11_n_0),
        .I2(g9314_INST_0_i_8_n_0),
        .I3(g614),
        .I4(g9280_INST_0_i_15_n_0),
        .I5(g9314_INST_0_i_9_n_0),
        .O(g9314_INST_0_i_3_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    g9314_INST_0_i_4
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9280_INST_0_i_19_n_0),
        .I2(g146),
        .O(g9314_INST_0_i_4_n_0));
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    g9314_INST_0_i_5
       (.I0(g9299_INST_0_i_4_n_0),
        .I1(g9314_INST_0_i_10_n_0),
        .I2(g9299_INST_0_i_14_n_0),
        .I3(g759),
        .I4(g9299_INST_0_i_15_n_0),
        .I5(g767),
        .O(g9314_INST_0_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF4F44FFFFFFFF)) 
    g9314_INST_0_i_6
       (.I0(g9299_INST_0_i_32_n_0),
        .I1(g751),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g498),
        .I4(g9314_INST_0_i_11_n_0),
        .I5(g9280_INST_0_i_6_n_0),
        .O(g9314_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9314_INST_0_i_7
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g563),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_25_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g601),
        .O(g9314_INST_0_i_7_n_0));
  LUT4 #(
    .INIT(16'hFEFF)) 
    g9314_INST_0_i_8
       (.I0(g9305_INST_0_i_6_n_0),
        .I1(g746_i_2_n_0),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g417),
        .O(g9314_INST_0_i_8_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9314_INST_0_i_9
       (.I0(g114),
        .I1(g9305_INST_0_i_6_n_0),
        .I2(g706_i_2_n_0),
        .I3(g9299_INST_0_i_16_n_0),
        .O(g9314_INST_0_i_9_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    g933_i_1
       (.I0(g933),
        .I1(g929),
        .O(g5166));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g933_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5166),
        .Q(g933));
  LUT3 #(
    .INIT(8'h8A)) 
    g936_i_1
       (.I0(g942),
        .I1(g936),
        .I2(g940),
        .O(g5168));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g936_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5168),
        .Q(g936));
  LUT6 #(
    .INIT(64'hE22E2EE2FFFFFFFF)) 
    g9378_INST_0
       (.I0(g7480),
        .I1(g44),
        .I2(g9378_INST_0_i_2_n_0),
        .I3(g9378_INST_0_i_3_n_0),
        .I4(g9378_INST_0_i_4_n_0),
        .I5(g62),
        .O(g9378));
  LUT5 #(
    .INIT(32'h4FB0B04F)) 
    g9378_INST_0_i_1
       (.I0(g45),
        .I1(g44),
        .I2(g47),
        .I3(g9378_INST_0_i_5_n_0),
        .I4(g9378_INST_0_i_6_n_0),
        .O(g7480));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    g9378_INST_0_i_10
       (.I0(g9299_INST_0_i_21_n_0),
        .I1(g9378_INST_0_i_23_n_0),
        .I2(g9280_INST_0_i_6_n_0),
        .I3(g9378_INST_0_i_24_n_0),
        .I4(g9378_INST_0_i_25_n_0),
        .I5(g9299_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    g9378_INST_0_i_11
       (.I0(g9378_INST_0_i_26_n_0),
        .I1(g300),
        .I2(g9378_INST_0_i_27_n_0),
        .I3(g348),
        .I4(g9310_INST_0_i_13_n_0),
        .O(g9378_INST_0_i_11_n_0));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    g9378_INST_0_i_12
       (.I0(g9297_INST_0_i_9_n_0),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g68),
        .I3(g610),
        .I4(g9280_INST_0_i_19_n_0),
        .I5(g154),
        .O(g9378_INST_0_i_12_n_0));
  LUT6 #(
    .INIT(64'h44444F4444444444)) 
    g9378_INST_0_i_13
       (.I0(g9280_INST_0_i_18_n_0),
        .I1(g130),
        .I2(g9297_INST_0_i_9_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g618),
        .O(g9378_INST_0_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    g9378_INST_0_i_14
       (.I0(g9305_INST_0_i_14_n_0),
        .I1(g9310_INST_0_i_9_n_0),
        .I2(g605),
        .I3(g9297_INST_0_i_17_n_0),
        .I4(g381),
        .I5(g9378_INST_0_i_28_n_0),
        .O(g9378_INST_0_i_14_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_15
       (.I0(g9378_INST_0_i_29_n_0),
        .I1(g597),
        .I2(g9297_INST_0_i_8_n_0),
        .I3(g219),
        .I4(g9305_INST_0_i_23_n_0),
        .O(g9378_INST_0_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    g9378_INST_0_i_16
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g74),
        .I3(g77),
        .I4(g71),
        .I5(g68),
        .O(g9378_INST_0_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    g9378_INST_0_i_17
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g9299_INST_0_i_17_n_0),
        .I2(g71),
        .I3(g74),
        .I4(g77),
        .I5(g68),
        .O(g9378_INST_0_i_17_n_0));
  LUT6 #(
    .INIT(64'hEFEEFFFFEFEEEFEE)) 
    g9378_INST_0_i_18
       (.I0(g9378_INST_0_i_30_n_0),
        .I1(g9378_INST_0_i_31_n_0),
        .I2(g4_i_3_n_0),
        .I3(g100),
        .I4(g9310_INST_0_i_9_n_0),
        .I5(g606),
        .O(g9378_INST_0_i_18_n_0));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    g9378_INST_0_i_19
       (.I0(g432),
        .I1(g9378_INST_0_i_32_n_0),
        .I2(g547),
        .I3(g9297_INST_0_i_11_n_0),
        .I4(g9310_INST_0_i_13_n_0),
        .I5(g351),
        .O(g9378_INST_0_i_19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g9378_INST_0_i_2
       (.I0(g9360),
        .I1(g9280_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    g9378_INST_0_i_20
       (.I0(g9297_INST_0_i_8_n_0),
        .I1(g598),
        .I2(g222),
        .I3(g9305_INST_0_i_23_n_0),
        .I4(g9378_INST_0_i_33_n_0),
        .O(g9378_INST_0_i_20_n_0));
  LUT5 #(
    .INIT(32'h10FF1010)) 
    g9378_INST_0_i_21
       (.I0(g7283_INST_0_i_2_n_0),
        .I1(g498_i_2_n_0),
        .I2(g630),
        .I3(g9299_INST_0_i_24_n_0),
        .I4(g270),
        .O(g9378_INST_0_i_21_n_0));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    g9378_INST_0_i_22
       (.I0(g9310_INST_0_i_14_n_0),
        .I1(g181),
        .I2(g134),
        .I3(g9280_INST_0_i_18_n_0),
        .I4(g158),
        .I5(g9280_INST_0_i_19_n_0),
        .O(g9378_INST_0_i_22_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_23
       (.I0(g9299_INST_0_i_18_n_0),
        .I1(g513),
        .I2(g9305_INST_0_i_30_n_0),
        .I3(g652),
        .I4(g9299_INST_0_i_20_n_0),
        .O(g9378_INST_0_i_23_n_0));
  LUT6 #(
    .INIT(64'h7707770700007707)) 
    g9378_INST_0_i_24
       (.I0(g9299_INST_0_i_11_n_0),
        .I1(g863),
        .I2(g2),
        .I3(g9378_INST_0_i_16_n_0),
        .I4(g846),
        .I5(g9378_INST_0_i_17_n_0),
        .O(g9378_INST_0_i_24_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    g9378_INST_0_i_25
       (.I0(g9312_INST_0_i_9_n_0),
        .I1(g772),
        .I2(g9299_INST_0_i_15_n_0),
        .I3(g764),
        .I4(g9299_INST_0_i_14_n_0),
        .O(g9378_INST_0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_26
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g68),
        .I2(g71),
        .I3(g77),
        .I4(g74),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_26_n_0));
  LUT6 #(
    .INIT(64'h0004000F00040004)) 
    g9378_INST_0_i_27
       (.I0(g9280_INST_0_i_35_n_0),
        .I1(g267),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9305_INST_0_i_6_n_0),
        .I4(g7283_INST_0_i_2_n_0),
        .I5(g180),
        .O(g9378_INST_0_i_27_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_28
       (.I0(g629),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g7283_INST_0_i_2_n_0),
        .O(g9378_INST_0_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_29
       (.I0(g9280_INST_0_i_34_n_0),
        .I1(g573),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g746_i_2_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g429),
        .O(g9378_INST_0_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAF355F3550C550C)) 
    g9378_INST_0_i_3
       (.I0(g9378_INST_0_i_7_n_0),
        .I1(g9305_INST_0_i_4_n_0),
        .I2(g9378_INST_0_i_8_n_0),
        .I3(g9299_INST_0_i_6_n_0),
        .I4(g9378_INST_0_i_9_n_0),
        .I5(g9378_INST_0_i_10_n_0),
        .O(g9378_INST_0_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000030200000002)) 
    g9378_INST_0_i_30
       (.I0(g611),
        .I1(g9308_INST_0_i_23_n_0),
        .I2(g9305_INST_0_i_6_n_0),
        .I3(g68),
        .I4(g9299_INST_0_i_16_n_0),
        .I5(g619),
        .O(g9378_INST_0_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000040F00000404)) 
    g9378_INST_0_i_31
       (.I0(g9280_INST_0_i_36_n_0),
        .I1(g303),
        .I2(g9299_INST_0_i_16_n_0),
        .I3(g9280_INST_0_i_31_n_0),
        .I4(g9305_INST_0_i_6_n_0),
        .I5(g384),
        .O(g9378_INST_0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    g9378_INST_0_i_32
       (.I0(g9299_INST_0_i_16_n_0),
        .I1(g74),
        .I2(g77),
        .I3(g71),
        .I4(g68),
        .I5(g9305_INST_0_i_6_n_0),
        .O(g9378_INST_0_i_32_n_0));
  LUT4 #(
    .INIT(16'h0002)) 
    g9378_INST_0_i_33
       (.I0(g622),
        .I1(g9299_INST_0_i_16_n_0),
        .I2(g9299_INST_0_i_17_n_0),
        .I3(g9305_INST_0_i_7_n_0),
        .O(g9378_INST_0_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_4
       (.I0(g9308_INST_0_i_1_n_0),
        .I1(g9376),
        .I2(g9312_INST_0_i_1_n_0),
        .I3(g9310_INST_0_i_1_n_0),
        .O(g9378_INST_0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_5
       (.I0(g4),
        .I1(g2),
        .I2(g3),
        .I3(g48),
        .O(g9378_INST_0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    g9378_INST_0_i_6
       (.I0(g8),
        .I1(g7),
        .I2(g6),
        .I3(g5),
        .O(g9378_INST_0_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_7
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_11_n_0),
        .I2(g9378_INST_0_i_12_n_0),
        .I3(g9378_INST_0_i_13_n_0),
        .I4(g9378_INST_0_i_14_n_0),
        .I5(g9378_INST_0_i_15_n_0),
        .O(g9378_INST_0_i_7_n_0));
  LUT6 #(
    .INIT(64'h000000000000D0DD)) 
    g9378_INST_0_i_8
       (.I0(g4),
        .I1(g9378_INST_0_i_16_n_0),
        .I2(g9378_INST_0_i_17_n_0),
        .I3(g843),
        .I4(g9305_INST_0_i_21_n_0),
        .I5(g9312_INST_0_i_9_n_0),
        .O(g9378_INST_0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g9378_INST_0_i_9
       (.I0(g9305_INST_0_i_1_n_0),
        .I1(g9378_INST_0_i_18_n_0),
        .I2(g9378_INST_0_i_19_n_0),
        .I3(g9378_INST_0_i_20_n_0),
        .I4(g9378_INST_0_i_21_n_0),
        .I5(g9378_INST_0_i_22_n_0),
        .O(g9378_INST_0_i_9_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g93_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g89),
        .Q(g93));
  LUT5 #(
    .INIT(32'h06666666)) 
    g940_i_1
       (.I0(g936),
        .I1(g940),
        .I2(g959),
        .I3(g955),
        .I4(g945),
        .O(g5735));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g940_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5735),
        .Q(g940));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g942_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g941),
        .Q(g942));
  LUT4 #(
    .INIT(16'hFB08)) 
    g943_i_1
       (.I0(g48),
        .I1(g936),
        .I2(g940),
        .I3(g954),
        .O(g8671));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g943_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8671),
        .Q(g943));
  LUT3 #(
    .INIT(8'h34)) 
    g944_i_1
       (.I0(g943),
        .I1(g940),
        .I2(g936),
        .O(g6372));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g944_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6372),
        .Q(g944));
  LUT3 #(
    .INIT(8'h6A)) 
    g945_i_1
       (.I0(g945),
        .I1(g955),
        .I2(g959),
        .O(g5170));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g945_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5170),
        .Q(g945));
  LUT3 #(
    .INIT(8'hEF)) 
    g948_i_1
       (.I0(g8),
        .I1(g940),
        .I2(g936),
        .O(g8664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g948_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8664),
        .Q(g948));
  LUT4 #(
    .INIT(16'hFB08)) 
    g949_i_1
       (.I0(g7),
        .I1(g936),
        .I2(g940),
        .I3(g948),
        .O(g8665));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g949_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8665),
        .Q(g949));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g94_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g4),
        .Q(g94));
  LUT4 #(
    .INIT(16'hFB08)) 
    g950_i_1
       (.I0(g6),
        .I1(g936),
        .I2(g940),
        .I3(g949),
        .O(g8666));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g950_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8666),
        .Q(g950));
  LUT4 #(
    .INIT(16'hFB08)) 
    g951_i_1
       (.I0(g5),
        .I1(g936),
        .I2(g940),
        .I3(g950),
        .O(g8667));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g951_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8667),
        .Q(g951));
  LUT4 #(
    .INIT(16'hFB08)) 
    g952_i_1
       (.I0(g4),
        .I1(g936),
        .I2(g940),
        .I3(g951),
        .O(g8668));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g952_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8668),
        .Q(g952));
  LUT4 #(
    .INIT(16'hFB08)) 
    g953_i_1
       (.I0(g2),
        .I1(g936),
        .I2(g940),
        .I3(g952),
        .O(g8669));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g953_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8669),
        .Q(g953));
  LUT4 #(
    .INIT(16'hFB08)) 
    g954_i_1
       (.I0(g3),
        .I1(g936),
        .I2(g940),
        .I3(g953),
        .O(g8670));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g954_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8670),
        .Q(g954));
  LUT1 #(
    .INIT(2'h1)) 
    g955_i_1
       (.I0(g955),
        .O(g1707));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g955_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1707),
        .Q(g955));
  LUT2 #(
    .INIT(4'h6)) 
    g959_i_1
       (.I0(g959),
        .I1(g955),
        .O(g5169));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g959_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g5169),
        .Q(g959));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g95_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g94),
        .Q(g95));
  LUT3 #(
    .INIT(8'h80)) 
    g963_i_1
       (.I0(g976),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7406));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g963_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7406),
        .Q(g963));
  LUT3 #(
    .INIT(8'h80)) 
    g966_i_1
       (.I0(g973),
        .I1(g7103_INST_0_i_1_n_0),
        .I2(g43),
        .O(g7566));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g966_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7566),
        .Q(g966));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g969_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g966),
        .Q(g969));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g970_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g963),
        .Q(g970));
  LUT1 #(
    .INIT(2'h1)) 
    g971_i_1
       (.I0(g1034),
        .O(g1789));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g971_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1789),
        .Q(g971));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g972_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g979),
        .Q(g972));
  LUT3 #(
    .INIT(8'h10)) 
    g973_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g973_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g973_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g973_i_1_n_0),
        .Q(g973));
  LUT3 #(
    .INIT(8'h40)) 
    g976_i_1
       (.I0(g7103_INST_0_i_1_n_0),
        .I1(g1),
        .I2(g43),
        .O(g976_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g976_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g976_i_1_n_0),
        .Q(g976));
  LUT3 #(
    .INIT(8'h08)) 
    g979_i_1
       (.I0(g984),
        .I1(g43),
        .I2(g979),
        .O(g6664));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g979_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g6664),
        .Q(g979));
  LUT2 #(
    .INIT(4'h2)) 
    g984_i_1
       (.I0(g7566),
        .I1(g979),
        .O(g9133));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g984_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9133),
        .Q(g984));
  LUT4 #(
    .INIT(16'h000D)) 
    g985_i_1
       (.I0(g995),
        .I1(g990),
        .I2(g985),
        .I3(g43),
        .O(g7515));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g985_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7515),
        .Q(g985));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g98_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g95),
        .Q(g98));
  LUT3 #(
    .INIT(8'h06)) 
    g990_i_1
       (.I0(g990),
        .I1(g985),
        .I2(g43),
        .O(g7516));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g990_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g7516),
        .Q(g990));
  LUT4 #(
    .INIT(16'h1540)) 
    g995_i_1
       (.I0(g43),
        .I1(g985),
        .I2(g990),
        .I3(g995),
        .O(g995_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g995_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g995_i_1_n_0),
        .Q(g995));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g998_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g1005),
        .Q(g998));
  LUT4 #(
    .INIT(16'h0020)) 
    g999_i_1
       (.I0(g1006_INST_0_i_1_n_0),
        .I1(g1000),
        .I2(g998),
        .I3(g1),
        .O(g8865));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g999_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g8865),
        .Q(g999));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  (* s = "true" *) 
  FDCE #(
    .INIT(1'b0)) 
    g99_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g2),
        .Q(g99));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* SHREG_EXTRACT = "no" *) 
  FDCE #(
    .INIT(1'b0)) 
    g9_reg
       (.C(blif_clk_net),
        .CE(1'b1),
        .CLR(blif_reset_net),
        .D(g9),
        .Q(g9));
endmodule
`ifndef GLBL
`define GLBL
`timescale  1 ps / 1 ps

module glbl ();

    parameter ROC_WIDTH = 100000;
    parameter TOC_WIDTH = 0;

//--------   STARTUP Globals --------------
    wire GSR;
    wire GTS;
    wire GWE;
    wire PRLD;
    tri1 p_up_tmp;
    tri (weak1, strong0) PLL_LOCKG = p_up_tmp;

    wire PROGB_GLBL;
    wire CCLKO_GLBL;
    wire FCSBO_GLBL;
    wire [3:0] DO_GLBL;
    wire [3:0] DI_GLBL;
   
    reg GSR_int;
    reg GTS_int;
    reg PRLD_int;

//--------   JTAG Globals --------------
    wire JTAG_TDO_GLBL;
    wire JTAG_TCK_GLBL;
    wire JTAG_TDI_GLBL;
    wire JTAG_TMS_GLBL;
    wire JTAG_TRST_GLBL;

    reg JTAG_CAPTURE_GLBL;
    reg JTAG_RESET_GLBL;
    reg JTAG_SHIFT_GLBL;
    reg JTAG_UPDATE_GLBL;
    reg JTAG_RUNTEST_GLBL;

    reg JTAG_SEL1_GLBL = 0;
    reg JTAG_SEL2_GLBL = 0 ;
    reg JTAG_SEL3_GLBL = 0;
    reg JTAG_SEL4_GLBL = 0;

    reg JTAG_USER_TDO1_GLBL = 1'bz;
    reg JTAG_USER_TDO2_GLBL = 1'bz;
    reg JTAG_USER_TDO3_GLBL = 1'bz;
    reg JTAG_USER_TDO4_GLBL = 1'bz;

    assign (strong1, weak0) GSR = GSR_int;
    assign (strong1, weak0) GTS = GTS_int;
    assign (weak1, weak0) PRLD = PRLD_int;

    initial begin
	GSR_int = 1'b1;
	PRLD_int = 1'b1;
	#(ROC_WIDTH)
	GSR_int = 1'b0;
	PRLD_int = 1'b0;
    end

    initial begin
	GTS_int = 1'b1;
	#(TOC_WIDTH)
	GTS_int = 1'b0;
    end

endmodule
`endif
