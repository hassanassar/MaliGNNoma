`timescale 1 ps / 1 ps
`define XIL_TIMING

module DSP48E2_UNIQ_BASE_
   (ACOUT,
    BCOUT,
    CARRYCASCOUT,
    CARRYOUT,
    MULTSIGNOUT,
    OVERFLOW,
    PATTERNBDETECT,
    PATTERNDETECT,
    PCOUT,
    P,
    UNDERFLOW,
    XOROUT,
    ACIN,
    ALUMODE,
    A,
    BCIN,
    B,
    CARRYCASCIN,
    CARRYIN,
    CARRYINSEL,
    CEA1,
    CEA2,
    CEAD,
    CEALUMODE,
    CEB1,
    CEB2,
    CEC,
    CECARRYIN,
    CECTRL,
    CED,
    CEINMODE,
    CEM,
    CEP,
    CLK,
    C,
    D,
    INMODE,
    MULTSIGNIN,
    OPMODE,
    PCIN,
    RSTA,
    RSTALLCARRYIN,
    RSTALUMODE,
    RSTB,
    RSTC,
    RSTCTRL,
    RSTD,
    RSTINMODE,
    RSTM,
    RSTP);
  output [29:0]ACOUT;
  output [17:0]BCOUT;
  output CARRYCASCOUT;
  output [3:0]CARRYOUT;
  output MULTSIGNOUT;
  output OVERFLOW;
  output PATTERNBDETECT;
  output PATTERNDETECT;
  output [47:0]PCOUT;
  output [47:0]P;
  output UNDERFLOW;
  output [7:0]XOROUT;
  input [29:0]ACIN;
  input [3:0]ALUMODE;
  input [29:0]A;
  input [17:0]BCIN;
  input [17:0]B;
  input CARRYCASCIN;
  input CARRYIN;
  input [2:0]CARRYINSEL;
  input CEA1;
  input CEA2;
  input CEAD;
  input CEALUMODE;
  input CEB1;
  input CEB2;
  input CEC;
  input CECARRYIN;
  input CECTRL;
  input CED;
  input CEINMODE;
  input CEM;
  input CEP;
  input CLK;
  input [47:0]C;
  input [26:0]D;
  input [4:0]INMODE;
  input MULTSIGNIN;
  input [8:0]OPMODE;
  input [47:0]PCIN;
  input RSTA;
  input RSTALLCARRYIN;
  input RSTALUMODE;
  input RSTB;
  input RSTC;
  input RSTCTRL;
  input RSTD;
  input RSTINMODE;
  input RSTM;
  input RSTP;

  wire \ACIN[0] ;
  wire \ACIN[10] ;
  wire \ACIN[11] ;
  wire \ACIN[12] ;
  wire \ACIN[13] ;
  wire \ACIN[14] ;
  wire \ACIN[15] ;
  wire \ACIN[16] ;
  wire \ACIN[17] ;
  wire \ACIN[18] ;
  wire \ACIN[19] ;
  wire \ACIN[1] ;
  wire \ACIN[20] ;
  wire \ACIN[21] ;
  wire \ACIN[22] ;
  wire \ACIN[23] ;
  wire \ACIN[24] ;
  wire \ACIN[25] ;
  wire \ACIN[26] ;
  wire \ACIN[27] ;
  wire \ACIN[28] ;
  wire \ACIN[29] ;
  wire \ACIN[2] ;
  wire \ACIN[3] ;
  wire \ACIN[4] ;
  wire \ACIN[5] ;
  wire \ACIN[6] ;
  wire \ACIN[7] ;
  wire \ACIN[8] ;
  wire \ACIN[9] ;
  wire \ACOUT[0] ;
  wire \ACOUT[10] ;
  wire \ACOUT[11] ;
  wire \ACOUT[12] ;
  wire \ACOUT[13] ;
  wire \ACOUT[14] ;
  wire \ACOUT[15] ;
  wire \ACOUT[16] ;
  wire \ACOUT[17] ;
  wire \ACOUT[18] ;
  wire \ACOUT[19] ;
  wire \ACOUT[1] ;
  wire \ACOUT[20] ;
  wire \ACOUT[21] ;
  wire \ACOUT[22] ;
  wire \ACOUT[23] ;
  wire \ACOUT[24] ;
  wire \ACOUT[25] ;
  wire \ACOUT[26] ;
  wire \ACOUT[27] ;
  wire \ACOUT[28] ;
  wire \ACOUT[29] ;
  wire \ACOUT[2] ;
  wire \ACOUT[3] ;
  wire \ACOUT[4] ;
  wire \ACOUT[5] ;
  wire \ACOUT[6] ;
  wire \ACOUT[7] ;
  wire \ACOUT[8] ;
  wire \ACOUT[9] ;
  wire \ALUMODE[0] ;
  wire \ALUMODE[1] ;
  wire \ALUMODE[2] ;
  wire \ALUMODE[3] ;
  wire \A[0] ;
  wire \A[10] ;
  wire \A[11] ;
  wire \A[12] ;
  wire \A[13] ;
  wire \A[14] ;
  wire \A[15] ;
  wire \A[16] ;
  wire \A[17] ;
  wire \A[18] ;
  wire \A[19] ;
  wire \A[1] ;
  wire \A[20] ;
  wire \A[21] ;
  wire \A[22] ;
  wire \A[23] ;
  wire \A[24] ;
  wire \A[25] ;
  wire \A[26] ;
  wire \A[27] ;
  wire \A[28] ;
  wire \A[29] ;
  wire \A[2] ;
  wire \A[3] ;
  wire \A[4] ;
  wire \A[5] ;
  wire \A[6] ;
  wire \A[7] ;
  wire \A[8] ;
  wire \A[9] ;
  wire \BCIN[0] ;
  wire \BCIN[10] ;
  wire \BCIN[11] ;
  wire \BCIN[12] ;
  wire \BCIN[13] ;
  wire \BCIN[14] ;
  wire \BCIN[15] ;
  wire \BCIN[16] ;
  wire \BCIN[17] ;
  wire \BCIN[1] ;
  wire \BCIN[2] ;
  wire \BCIN[3] ;
  wire \BCIN[4] ;
  wire \BCIN[5] ;
  wire \BCIN[6] ;
  wire \BCIN[7] ;
  wire \BCIN[8] ;
  wire \BCIN[9] ;
  wire \BCOUT[0] ;
  wire \BCOUT[10] ;
  wire \BCOUT[11] ;
  wire \BCOUT[12] ;
  wire \BCOUT[13] ;
  wire \BCOUT[14] ;
  wire \BCOUT[15] ;
  wire \BCOUT[16] ;
  wire \BCOUT[17] ;
  wire \BCOUT[1] ;
  wire \BCOUT[2] ;
  wire \BCOUT[3] ;
  wire \BCOUT[4] ;
  wire \BCOUT[5] ;
  wire \BCOUT[6] ;
  wire \BCOUT[7] ;
  wire \BCOUT[8] ;
  wire \BCOUT[9] ;
  wire \B[0] ;
  wire \B[10] ;
  wire \B[11] ;
  wire \B[12] ;
  wire \B[13] ;
  wire \B[14] ;
  wire \B[15] ;
  wire \B[16] ;
  wire \B[17] ;
  wire \B[1] ;
  wire \B[2] ;
  wire \B[3] ;
  wire \B[4] ;
  wire \B[5] ;
  wire \B[6] ;
  wire \B[7] ;
  wire \B[8] ;
  wire \B[9] ;
  wire CARRYCASCIN;
  wire CARRYCASCOUT;
  wire CARRYIN;
  wire \CARRYINSEL[0] ;
  wire \CARRYINSEL[1] ;
  wire \CARRYINSEL[2] ;
  wire \CARRYOUT[0] ;
  wire \CARRYOUT[1] ;
  wire \CARRYOUT[2] ;
  wire \CARRYOUT[3] ;
  wire CEA1;
  wire CEA2;
  wire CEAD;
  wire CEALUMODE;
  wire CEB1;
  wire CEB2;
  wire CEC;
  wire CECARRYIN;
  wire CECTRL;
  wire CED;
  wire CEINMODE;
  wire CEM;
  wire CEP;
  wire CLK;
  wire \C[0] ;
  wire \C[10] ;
  wire \C[11] ;
  wire \C[12] ;
  wire \C[13] ;
  wire \C[14] ;
  wire \C[15] ;
  wire \C[16] ;
  wire \C[17] ;
  wire \C[18] ;
  wire \C[19] ;
  wire \C[1] ;
  wire \C[20] ;
  wire \C[21] ;
  wire \C[22] ;
  wire \C[23] ;
  wire \C[24] ;
  wire \C[25] ;
  wire \C[26] ;
  wire \C[27] ;
  wire \C[28] ;
  wire \C[29] ;
  wire \C[2] ;
  wire \C[30] ;
  wire \C[31] ;
  wire \C[32] ;
  wire \C[33] ;
  wire \C[34] ;
  wire \C[35] ;
  wire \C[36] ;
  wire \C[37] ;
  wire \C[38] ;
  wire \C[39] ;
  wire \C[3] ;
  wire \C[40] ;
  wire \C[41] ;
  wire \C[42] ;
  wire \C[43] ;
  wire \C[44] ;
  wire \C[45] ;
  wire \C[46] ;
  wire \C[47] ;
  wire \C[4] ;
  wire \C[5] ;
  wire \C[6] ;
  wire \C[7] ;
  wire \C[8] ;
  wire \C[9] ;
  wire \DSP_ALU.ALUMODE10 ;
  wire \DSP_ALU.ALU_OUT<0> ;
  wire \DSP_ALU.ALU_OUT<10> ;
  wire \DSP_ALU.ALU_OUT<11> ;
  wire \DSP_ALU.ALU_OUT<12> ;
  wire \DSP_ALU.ALU_OUT<13> ;
  wire \DSP_ALU.ALU_OUT<14> ;
  wire \DSP_ALU.ALU_OUT<15> ;
  wire \DSP_ALU.ALU_OUT<16> ;
  wire \DSP_ALU.ALU_OUT<17> ;
  wire \DSP_ALU.ALU_OUT<18> ;
  wire \DSP_ALU.ALU_OUT<19> ;
  wire \DSP_ALU.ALU_OUT<1> ;
  wire \DSP_ALU.ALU_OUT<20> ;
  wire \DSP_ALU.ALU_OUT<21> ;
  wire \DSP_ALU.ALU_OUT<22> ;
  wire \DSP_ALU.ALU_OUT<23> ;
  wire \DSP_ALU.ALU_OUT<24> ;
  wire \DSP_ALU.ALU_OUT<25> ;
  wire \DSP_ALU.ALU_OUT<26> ;
  wire \DSP_ALU.ALU_OUT<27> ;
  wire \DSP_ALU.ALU_OUT<28> ;
  wire \DSP_ALU.ALU_OUT<29> ;
  wire \DSP_ALU.ALU_OUT<2> ;
  wire \DSP_ALU.ALU_OUT<30> ;
  wire \DSP_ALU.ALU_OUT<31> ;
  wire \DSP_ALU.ALU_OUT<32> ;
  wire \DSP_ALU.ALU_OUT<33> ;
  wire \DSP_ALU.ALU_OUT<34> ;
  wire \DSP_ALU.ALU_OUT<35> ;
  wire \DSP_ALU.ALU_OUT<36> ;
  wire \DSP_ALU.ALU_OUT<37> ;
  wire \DSP_ALU.ALU_OUT<38> ;
  wire \DSP_ALU.ALU_OUT<39> ;
  wire \DSP_ALU.ALU_OUT<3> ;
  wire \DSP_ALU.ALU_OUT<40> ;
  wire \DSP_ALU.ALU_OUT<41> ;
  wire \DSP_ALU.ALU_OUT<42> ;
  wire \DSP_ALU.ALU_OUT<43> ;
  wire \DSP_ALU.ALU_OUT<44> ;
  wire \DSP_ALU.ALU_OUT<45> ;
  wire \DSP_ALU.ALU_OUT<46> ;
  wire \DSP_ALU.ALU_OUT<47> ;
  wire \DSP_ALU.ALU_OUT<4> ;
  wire \DSP_ALU.ALU_OUT<5> ;
  wire \DSP_ALU.ALU_OUT<6> ;
  wire \DSP_ALU.ALU_OUT<7> ;
  wire \DSP_ALU.ALU_OUT<8> ;
  wire \DSP_ALU.ALU_OUT<9> ;
  wire \DSP_ALU.COUT<0> ;
  wire \DSP_ALU.COUT<1> ;
  wire \DSP_ALU.COUT<2> ;
  wire \DSP_ALU.COUT<3> ;
  wire \DSP_ALU.MULTSIGN_ALU ;
  wire \DSP_ALU.XOR_MX<0> ;
  wire \DSP_ALU.XOR_MX<1> ;
  wire \DSP_ALU.XOR_MX<2> ;
  wire \DSP_ALU.XOR_MX<3> ;
  wire \DSP_ALU.XOR_MX<4> ;
  wire \DSP_ALU.XOR_MX<5> ;
  wire \DSP_ALU.XOR_MX<6> ;
  wire \DSP_ALU.XOR_MX<7> ;
  wire \DSP_A_B_DATA.A1_DATA<0> ;
  wire \DSP_A_B_DATA.A1_DATA<10> ;
  wire \DSP_A_B_DATA.A1_DATA<11> ;
  wire \DSP_A_B_DATA.A1_DATA<12> ;
  wire \DSP_A_B_DATA.A1_DATA<13> ;
  wire \DSP_A_B_DATA.A1_DATA<14> ;
  wire \DSP_A_B_DATA.A1_DATA<15> ;
  wire \DSP_A_B_DATA.A1_DATA<16> ;
  wire \DSP_A_B_DATA.A1_DATA<17> ;
  wire \DSP_A_B_DATA.A1_DATA<18> ;
  wire \DSP_A_B_DATA.A1_DATA<19> ;
  wire \DSP_A_B_DATA.A1_DATA<1> ;
  wire \DSP_A_B_DATA.A1_DATA<20> ;
  wire \DSP_A_B_DATA.A1_DATA<21> ;
  wire \DSP_A_B_DATA.A1_DATA<22> ;
  wire \DSP_A_B_DATA.A1_DATA<23> ;
  wire \DSP_A_B_DATA.A1_DATA<24> ;
  wire \DSP_A_B_DATA.A1_DATA<25> ;
  wire \DSP_A_B_DATA.A1_DATA<26> ;
  wire \DSP_A_B_DATA.A1_DATA<2> ;
  wire \DSP_A_B_DATA.A1_DATA<3> ;
  wire \DSP_A_B_DATA.A1_DATA<4> ;
  wire \DSP_A_B_DATA.A1_DATA<5> ;
  wire \DSP_A_B_DATA.A1_DATA<6> ;
  wire \DSP_A_B_DATA.A1_DATA<7> ;
  wire \DSP_A_B_DATA.A1_DATA<8> ;
  wire \DSP_A_B_DATA.A1_DATA<9> ;
  wire \DSP_A_B_DATA.A2_DATA<0> ;
  wire \DSP_A_B_DATA.A2_DATA<10> ;
  wire \DSP_A_B_DATA.A2_DATA<11> ;
  wire \DSP_A_B_DATA.A2_DATA<12> ;
  wire \DSP_A_B_DATA.A2_DATA<13> ;
  wire \DSP_A_B_DATA.A2_DATA<14> ;
  wire \DSP_A_B_DATA.A2_DATA<15> ;
  wire \DSP_A_B_DATA.A2_DATA<16> ;
  wire \DSP_A_B_DATA.A2_DATA<17> ;
  wire \DSP_A_B_DATA.A2_DATA<18> ;
  wire \DSP_A_B_DATA.A2_DATA<19> ;
  wire \DSP_A_B_DATA.A2_DATA<1> ;
  wire \DSP_A_B_DATA.A2_DATA<20> ;
  wire \DSP_A_B_DATA.A2_DATA<21> ;
  wire \DSP_A_B_DATA.A2_DATA<22> ;
  wire \DSP_A_B_DATA.A2_DATA<23> ;
  wire \DSP_A_B_DATA.A2_DATA<24> ;
  wire \DSP_A_B_DATA.A2_DATA<25> ;
  wire \DSP_A_B_DATA.A2_DATA<26> ;
  wire \DSP_A_B_DATA.A2_DATA<2> ;
  wire \DSP_A_B_DATA.A2_DATA<3> ;
  wire \DSP_A_B_DATA.A2_DATA<4> ;
  wire \DSP_A_B_DATA.A2_DATA<5> ;
  wire \DSP_A_B_DATA.A2_DATA<6> ;
  wire \DSP_A_B_DATA.A2_DATA<7> ;
  wire \DSP_A_B_DATA.A2_DATA<8> ;
  wire \DSP_A_B_DATA.A2_DATA<9> ;
  wire \DSP_A_B_DATA.A_ALU<0> ;
  wire \DSP_A_B_DATA.A_ALU<10> ;
  wire \DSP_A_B_DATA.A_ALU<11> ;
  wire \DSP_A_B_DATA.A_ALU<12> ;
  wire \DSP_A_B_DATA.A_ALU<13> ;
  wire \DSP_A_B_DATA.A_ALU<14> ;
  wire \DSP_A_B_DATA.A_ALU<15> ;
  wire \DSP_A_B_DATA.A_ALU<16> ;
  wire \DSP_A_B_DATA.A_ALU<17> ;
  wire \DSP_A_B_DATA.A_ALU<18> ;
  wire \DSP_A_B_DATA.A_ALU<19> ;
  wire \DSP_A_B_DATA.A_ALU<1> ;
  wire \DSP_A_B_DATA.A_ALU<20> ;
  wire \DSP_A_B_DATA.A_ALU<21> ;
  wire \DSP_A_B_DATA.A_ALU<22> ;
  wire \DSP_A_B_DATA.A_ALU<23> ;
  wire \DSP_A_B_DATA.A_ALU<24> ;
  wire \DSP_A_B_DATA.A_ALU<25> ;
  wire \DSP_A_B_DATA.A_ALU<26> ;
  wire \DSP_A_B_DATA.A_ALU<27> ;
  wire \DSP_A_B_DATA.A_ALU<28> ;
  wire \DSP_A_B_DATA.A_ALU<29> ;
  wire \DSP_A_B_DATA.A_ALU<2> ;
  wire \DSP_A_B_DATA.A_ALU<3> ;
  wire \DSP_A_B_DATA.A_ALU<4> ;
  wire \DSP_A_B_DATA.A_ALU<5> ;
  wire \DSP_A_B_DATA.A_ALU<6> ;
  wire \DSP_A_B_DATA.A_ALU<7> ;
  wire \DSP_A_B_DATA.A_ALU<8> ;
  wire \DSP_A_B_DATA.A_ALU<9> ;
  wire \DSP_A_B_DATA.B1_DATA<0> ;
  wire \DSP_A_B_DATA.B1_DATA<10> ;
  wire \DSP_A_B_DATA.B1_DATA<11> ;
  wire \DSP_A_B_DATA.B1_DATA<12> ;
  wire \DSP_A_B_DATA.B1_DATA<13> ;
  wire \DSP_A_B_DATA.B1_DATA<14> ;
  wire \DSP_A_B_DATA.B1_DATA<15> ;
  wire \DSP_A_B_DATA.B1_DATA<16> ;
  wire \DSP_A_B_DATA.B1_DATA<17> ;
  wire \DSP_A_B_DATA.B1_DATA<1> ;
  wire \DSP_A_B_DATA.B1_DATA<2> ;
  wire \DSP_A_B_DATA.B1_DATA<3> ;
  wire \DSP_A_B_DATA.B1_DATA<4> ;
  wire \DSP_A_B_DATA.B1_DATA<5> ;
  wire \DSP_A_B_DATA.B1_DATA<6> ;
  wire \DSP_A_B_DATA.B1_DATA<7> ;
  wire \DSP_A_B_DATA.B1_DATA<8> ;
  wire \DSP_A_B_DATA.B1_DATA<9> ;
  wire \DSP_A_B_DATA.B2_DATA<0> ;
  wire \DSP_A_B_DATA.B2_DATA<10> ;
  wire \DSP_A_B_DATA.B2_DATA<11> ;
  wire \DSP_A_B_DATA.B2_DATA<12> ;
  wire \DSP_A_B_DATA.B2_DATA<13> ;
  wire \DSP_A_B_DATA.B2_DATA<14> ;
  wire \DSP_A_B_DATA.B2_DATA<15> ;
  wire \DSP_A_B_DATA.B2_DATA<16> ;
  wire \DSP_A_B_DATA.B2_DATA<17> ;
  wire \DSP_A_B_DATA.B2_DATA<1> ;
  wire \DSP_A_B_DATA.B2_DATA<2> ;
  wire \DSP_A_B_DATA.B2_DATA<3> ;
  wire \DSP_A_B_DATA.B2_DATA<4> ;
  wire \DSP_A_B_DATA.B2_DATA<5> ;
  wire \DSP_A_B_DATA.B2_DATA<6> ;
  wire \DSP_A_B_DATA.B2_DATA<7> ;
  wire \DSP_A_B_DATA.B2_DATA<8> ;
  wire \DSP_A_B_DATA.B2_DATA<9> ;
  wire \DSP_A_B_DATA.B_ALU<0> ;
  wire \DSP_A_B_DATA.B_ALU<10> ;
  wire \DSP_A_B_DATA.B_ALU<11> ;
  wire \DSP_A_B_DATA.B_ALU<12> ;
  wire \DSP_A_B_DATA.B_ALU<13> ;
  wire \DSP_A_B_DATA.B_ALU<14> ;
  wire \DSP_A_B_DATA.B_ALU<15> ;
  wire \DSP_A_B_DATA.B_ALU<16> ;
  wire \DSP_A_B_DATA.B_ALU<17> ;
  wire \DSP_A_B_DATA.B_ALU<1> ;
  wire \DSP_A_B_DATA.B_ALU<2> ;
  wire \DSP_A_B_DATA.B_ALU<3> ;
  wire \DSP_A_B_DATA.B_ALU<4> ;
  wire \DSP_A_B_DATA.B_ALU<5> ;
  wire \DSP_A_B_DATA.B_ALU<6> ;
  wire \DSP_A_B_DATA.B_ALU<7> ;
  wire \DSP_A_B_DATA.B_ALU<8> ;
  wire \DSP_A_B_DATA.B_ALU<9> ;
  wire \DSP_C_DATA.C_DATA<0> ;
  wire \DSP_C_DATA.C_DATA<10> ;
  wire \DSP_C_DATA.C_DATA<11> ;
  wire \DSP_C_DATA.C_DATA<12> ;
  wire \DSP_C_DATA.C_DATA<13> ;
  wire \DSP_C_DATA.C_DATA<14> ;
  wire \DSP_C_DATA.C_DATA<15> ;
  wire \DSP_C_DATA.C_DATA<16> ;
  wire \DSP_C_DATA.C_DATA<17> ;
  wire \DSP_C_DATA.C_DATA<18> ;
  wire \DSP_C_DATA.C_DATA<19> ;
  wire \DSP_C_DATA.C_DATA<1> ;
  wire \DSP_C_DATA.C_DATA<20> ;
  wire \DSP_C_DATA.C_DATA<21> ;
  wire \DSP_C_DATA.C_DATA<22> ;
  wire \DSP_C_DATA.C_DATA<23> ;
  wire \DSP_C_DATA.C_DATA<24> ;
  wire \DSP_C_DATA.C_DATA<25> ;
  wire \DSP_C_DATA.C_DATA<26> ;
  wire \DSP_C_DATA.C_DATA<27> ;
  wire \DSP_C_DATA.C_DATA<28> ;
  wire \DSP_C_DATA.C_DATA<29> ;
  wire \DSP_C_DATA.C_DATA<2> ;
  wire \DSP_C_DATA.C_DATA<30> ;
  wire \DSP_C_DATA.C_DATA<31> ;
  wire \DSP_C_DATA.C_DATA<32> ;
  wire \DSP_C_DATA.C_DATA<33> ;
  wire \DSP_C_DATA.C_DATA<34> ;
  wire \DSP_C_DATA.C_DATA<35> ;
  wire \DSP_C_DATA.C_DATA<36> ;
  wire \DSP_C_DATA.C_DATA<37> ;
  wire \DSP_C_DATA.C_DATA<38> ;
  wire \DSP_C_DATA.C_DATA<39> ;
  wire \DSP_C_DATA.C_DATA<3> ;
  wire \DSP_C_DATA.C_DATA<40> ;
  wire \DSP_C_DATA.C_DATA<41> ;
  wire \DSP_C_DATA.C_DATA<42> ;
  wire \DSP_C_DATA.C_DATA<43> ;
  wire \DSP_C_DATA.C_DATA<44> ;
  wire \DSP_C_DATA.C_DATA<45> ;
  wire \DSP_C_DATA.C_DATA<46> ;
  wire \DSP_C_DATA.C_DATA<47> ;
  wire \DSP_C_DATA.C_DATA<4> ;
  wire \DSP_C_DATA.C_DATA<5> ;
  wire \DSP_C_DATA.C_DATA<6> ;
  wire \DSP_C_DATA.C_DATA<7> ;
  wire \DSP_C_DATA.C_DATA<8> ;
  wire \DSP_C_DATA.C_DATA<9> ;
  wire \DSP_MULTIPLIER.AMULT26 ;
  wire \DSP_MULTIPLIER.BMULT17 ;
  wire \DSP_MULTIPLIER.U<0> ;
  wire \DSP_MULTIPLIER.U<10> ;
  wire \DSP_MULTIPLIER.U<11> ;
  wire \DSP_MULTIPLIER.U<12> ;
  wire \DSP_MULTIPLIER.U<13> ;
  wire \DSP_MULTIPLIER.U<14> ;
  wire \DSP_MULTIPLIER.U<15> ;
  wire \DSP_MULTIPLIER.U<16> ;
  wire \DSP_MULTIPLIER.U<17> ;
  wire \DSP_MULTIPLIER.U<18> ;
  wire \DSP_MULTIPLIER.U<19> ;
  wire \DSP_MULTIPLIER.U<1> ;
  wire \DSP_MULTIPLIER.U<20> ;
  wire \DSP_MULTIPLIER.U<21> ;
  wire \DSP_MULTIPLIER.U<22> ;
  wire \DSP_MULTIPLIER.U<23> ;
  wire \DSP_MULTIPLIER.U<24> ;
  wire \DSP_MULTIPLIER.U<25> ;
  wire \DSP_MULTIPLIER.U<26> ;
  wire \DSP_MULTIPLIER.U<27> ;
  wire \DSP_MULTIPLIER.U<28> ;
  wire \DSP_MULTIPLIER.U<29> ;
  wire \DSP_MULTIPLIER.U<2> ;
  wire \DSP_MULTIPLIER.U<30> ;
  wire \DSP_MULTIPLIER.U<31> ;
  wire \DSP_MULTIPLIER.U<32> ;
  wire \DSP_MULTIPLIER.U<33> ;
  wire \DSP_MULTIPLIER.U<34> ;
  wire \DSP_MULTIPLIER.U<35> ;
  wire \DSP_MULTIPLIER.U<36> ;
  wire \DSP_MULTIPLIER.U<37> ;
  wire \DSP_MULTIPLIER.U<38> ;
  wire \DSP_MULTIPLIER.U<39> ;
  wire \DSP_MULTIPLIER.U<3> ;
  wire \DSP_MULTIPLIER.U<40> ;
  wire \DSP_MULTIPLIER.U<41> ;
  wire \DSP_MULTIPLIER.U<42> ;
  wire \DSP_MULTIPLIER.U<43> ;
  wire \DSP_MULTIPLIER.U<44> ;
  wire \DSP_MULTIPLIER.U<4> ;
  wire \DSP_MULTIPLIER.U<5> ;
  wire \DSP_MULTIPLIER.U<6> ;
  wire \DSP_MULTIPLIER.U<7> ;
  wire \DSP_MULTIPLIER.U<8> ;
  wire \DSP_MULTIPLIER.U<9> ;
  wire \DSP_MULTIPLIER.V<0> ;
  wire \DSP_MULTIPLIER.V<10> ;
  wire \DSP_MULTIPLIER.V<11> ;
  wire \DSP_MULTIPLIER.V<12> ;
  wire \DSP_MULTIPLIER.V<13> ;
  wire \DSP_MULTIPLIER.V<14> ;
  wire \DSP_MULTIPLIER.V<15> ;
  wire \DSP_MULTIPLIER.V<16> ;
  wire \DSP_MULTIPLIER.V<17> ;
  wire \DSP_MULTIPLIER.V<18> ;
  wire \DSP_MULTIPLIER.V<19> ;
  wire \DSP_MULTIPLIER.V<1> ;
  wire \DSP_MULTIPLIER.V<20> ;
  wire \DSP_MULTIPLIER.V<21> ;
  wire \DSP_MULTIPLIER.V<22> ;
  wire \DSP_MULTIPLIER.V<23> ;
  wire \DSP_MULTIPLIER.V<24> ;
  wire \DSP_MULTIPLIER.V<25> ;
  wire \DSP_MULTIPLIER.V<26> ;
  wire \DSP_MULTIPLIER.V<27> ;
  wire \DSP_MULTIPLIER.V<28> ;
  wire \DSP_MULTIPLIER.V<29> ;
  wire \DSP_MULTIPLIER.V<2> ;
  wire \DSP_MULTIPLIER.V<30> ;
  wire \DSP_MULTIPLIER.V<31> ;
  wire \DSP_MULTIPLIER.V<32> ;
  wire \DSP_MULTIPLIER.V<33> ;
  wire \DSP_MULTIPLIER.V<34> ;
  wire \DSP_MULTIPLIER.V<35> ;
  wire \DSP_MULTIPLIER.V<36> ;
  wire \DSP_MULTIPLIER.V<37> ;
  wire \DSP_MULTIPLIER.V<38> ;
  wire \DSP_MULTIPLIER.V<39> ;
  wire \DSP_MULTIPLIER.V<3> ;
  wire \DSP_MULTIPLIER.V<40> ;
  wire \DSP_MULTIPLIER.V<41> ;
  wire \DSP_MULTIPLIER.V<42> ;
  wire \DSP_MULTIPLIER.V<43> ;
  wire \DSP_MULTIPLIER.V<44> ;
  wire \DSP_MULTIPLIER.V<4> ;
  wire \DSP_MULTIPLIER.V<5> ;
  wire \DSP_MULTIPLIER.V<6> ;
  wire \DSP_MULTIPLIER.V<7> ;
  wire \DSP_MULTIPLIER.V<8> ;
  wire \DSP_MULTIPLIER.V<9> ;
  wire \DSP_M_DATA.U_DATA<0> ;
  wire \DSP_M_DATA.U_DATA<10> ;
  wire \DSP_M_DATA.U_DATA<11> ;
  wire \DSP_M_DATA.U_DATA<12> ;
  wire \DSP_M_DATA.U_DATA<13> ;
  wire \DSP_M_DATA.U_DATA<14> ;
  wire \DSP_M_DATA.U_DATA<15> ;
  wire \DSP_M_DATA.U_DATA<16> ;
  wire \DSP_M_DATA.U_DATA<17> ;
  wire \DSP_M_DATA.U_DATA<18> ;
  wire \DSP_M_DATA.U_DATA<19> ;
  wire \DSP_M_DATA.U_DATA<1> ;
  wire \DSP_M_DATA.U_DATA<20> ;
  wire \DSP_M_DATA.U_DATA<21> ;
  wire \DSP_M_DATA.U_DATA<22> ;
  wire \DSP_M_DATA.U_DATA<23> ;
  wire \DSP_M_DATA.U_DATA<24> ;
  wire \DSP_M_DATA.U_DATA<25> ;
  wire \DSP_M_DATA.U_DATA<26> ;
  wire \DSP_M_DATA.U_DATA<27> ;
  wire \DSP_M_DATA.U_DATA<28> ;
  wire \DSP_M_DATA.U_DATA<29> ;
  wire \DSP_M_DATA.U_DATA<2> ;
  wire \DSP_M_DATA.U_DATA<30> ;
  wire \DSP_M_DATA.U_DATA<31> ;
  wire \DSP_M_DATA.U_DATA<32> ;
  wire \DSP_M_DATA.U_DATA<33> ;
  wire \DSP_M_DATA.U_DATA<34> ;
  wire \DSP_M_DATA.U_DATA<35> ;
  wire \DSP_M_DATA.U_DATA<36> ;
  wire \DSP_M_DATA.U_DATA<37> ;
  wire \DSP_M_DATA.U_DATA<38> ;
  wire \DSP_M_DATA.U_DATA<39> ;
  wire \DSP_M_DATA.U_DATA<3> ;
  wire \DSP_M_DATA.U_DATA<40> ;
  wire \DSP_M_DATA.U_DATA<41> ;
  wire \DSP_M_DATA.U_DATA<42> ;
  wire \DSP_M_DATA.U_DATA<43> ;
  wire \DSP_M_DATA.U_DATA<44> ;
  wire \DSP_M_DATA.U_DATA<4> ;
  wire \DSP_M_DATA.U_DATA<5> ;
  wire \DSP_M_DATA.U_DATA<6> ;
  wire \DSP_M_DATA.U_DATA<7> ;
  wire \DSP_M_DATA.U_DATA<8> ;
  wire \DSP_M_DATA.U_DATA<9> ;
  wire \DSP_M_DATA.V_DATA<0> ;
  wire \DSP_M_DATA.V_DATA<10> ;
  wire \DSP_M_DATA.V_DATA<11> ;
  wire \DSP_M_DATA.V_DATA<12> ;
  wire \DSP_M_DATA.V_DATA<13> ;
  wire \DSP_M_DATA.V_DATA<14> ;
  wire \DSP_M_DATA.V_DATA<15> ;
  wire \DSP_M_DATA.V_DATA<16> ;
  wire \DSP_M_DATA.V_DATA<17> ;
  wire \DSP_M_DATA.V_DATA<18> ;
  wire \DSP_M_DATA.V_DATA<19> ;
  wire \DSP_M_DATA.V_DATA<1> ;
  wire \DSP_M_DATA.V_DATA<20> ;
  wire \DSP_M_DATA.V_DATA<21> ;
  wire \DSP_M_DATA.V_DATA<22> ;
  wire \DSP_M_DATA.V_DATA<23> ;
  wire \DSP_M_DATA.V_DATA<24> ;
  wire \DSP_M_DATA.V_DATA<25> ;
  wire \DSP_M_DATA.V_DATA<26> ;
  wire \DSP_M_DATA.V_DATA<27> ;
  wire \DSP_M_DATA.V_DATA<28> ;
  wire \DSP_M_DATA.V_DATA<29> ;
  wire \DSP_M_DATA.V_DATA<2> ;
  wire \DSP_M_DATA.V_DATA<30> ;
  wire \DSP_M_DATA.V_DATA<31> ;
  wire \DSP_M_DATA.V_DATA<32> ;
  wire \DSP_M_DATA.V_DATA<33> ;
  wire \DSP_M_DATA.V_DATA<34> ;
  wire \DSP_M_DATA.V_DATA<35> ;
  wire \DSP_M_DATA.V_DATA<36> ;
  wire \DSP_M_DATA.V_DATA<37> ;
  wire \DSP_M_DATA.V_DATA<38> ;
  wire \DSP_M_DATA.V_DATA<39> ;
  wire \DSP_M_DATA.V_DATA<3> ;
  wire \DSP_M_DATA.V_DATA<40> ;
  wire \DSP_M_DATA.V_DATA<41> ;
  wire \DSP_M_DATA.V_DATA<42> ;
  wire \DSP_M_DATA.V_DATA<43> ;
  wire \DSP_M_DATA.V_DATA<44> ;
  wire \DSP_M_DATA.V_DATA<4> ;
  wire \DSP_M_DATA.V_DATA<5> ;
  wire \DSP_M_DATA.V_DATA<6> ;
  wire \DSP_M_DATA.V_DATA<7> ;
  wire \DSP_M_DATA.V_DATA<8> ;
  wire \DSP_M_DATA.V_DATA<9> ;
  wire \DSP_OUTPUT.CCOUT_FB ;
  wire \DSP_OUTPUT.P_FDBK<0> ;
  wire \DSP_OUTPUT.P_FDBK<10> ;
  wire \DSP_OUTPUT.P_FDBK<11> ;
  wire \DSP_OUTPUT.P_FDBK<12> ;
  wire \DSP_OUTPUT.P_FDBK<13> ;
  wire \DSP_OUTPUT.P_FDBK<14> ;
  wire \DSP_OUTPUT.P_FDBK<15> ;
  wire \DSP_OUTPUT.P_FDBK<16> ;
  wire \DSP_OUTPUT.P_FDBK<17> ;
  wire \DSP_OUTPUT.P_FDBK<18> ;
  wire \DSP_OUTPUT.P_FDBK<19> ;
  wire \DSP_OUTPUT.P_FDBK<1> ;
  wire \DSP_OUTPUT.P_FDBK<20> ;
  wire \DSP_OUTPUT.P_FDBK<21> ;
  wire \DSP_OUTPUT.P_FDBK<22> ;
  wire \DSP_OUTPUT.P_FDBK<23> ;
  wire \DSP_OUTPUT.P_FDBK<24> ;
  wire \DSP_OUTPUT.P_FDBK<25> ;
  wire \DSP_OUTPUT.P_FDBK<26> ;
  wire \DSP_OUTPUT.P_FDBK<27> ;
  wire \DSP_OUTPUT.P_FDBK<28> ;
  wire \DSP_OUTPUT.P_FDBK<29> ;
  wire \DSP_OUTPUT.P_FDBK<2> ;
  wire \DSP_OUTPUT.P_FDBK<30> ;
  wire \DSP_OUTPUT.P_FDBK<31> ;
  wire \DSP_OUTPUT.P_FDBK<32> ;
  wire \DSP_OUTPUT.P_FDBK<33> ;
  wire \DSP_OUTPUT.P_FDBK<34> ;
  wire \DSP_OUTPUT.P_FDBK<35> ;
  wire \DSP_OUTPUT.P_FDBK<36> ;
  wire \DSP_OUTPUT.P_FDBK<37> ;
  wire \DSP_OUTPUT.P_FDBK<38> ;
  wire \DSP_OUTPUT.P_FDBK<39> ;
  wire \DSP_OUTPUT.P_FDBK<3> ;
  wire \DSP_OUTPUT.P_FDBK<40> ;
  wire \DSP_OUTPUT.P_FDBK<41> ;
  wire \DSP_OUTPUT.P_FDBK<42> ;
  wire \DSP_OUTPUT.P_FDBK<43> ;
  wire \DSP_OUTPUT.P_FDBK<44> ;
  wire \DSP_OUTPUT.P_FDBK<45> ;
  wire \DSP_OUTPUT.P_FDBK<46> ;
  wire \DSP_OUTPUT.P_FDBK<47> ;
  wire \DSP_OUTPUT.P_FDBK<4> ;
  wire \DSP_OUTPUT.P_FDBK<5> ;
  wire \DSP_OUTPUT.P_FDBK<6> ;
  wire \DSP_OUTPUT.P_FDBK<7> ;
  wire \DSP_OUTPUT.P_FDBK<8> ;
  wire \DSP_OUTPUT.P_FDBK<9> ;
  wire \DSP_OUTPUT.P_FDBK_47 ;
  wire \DSP_PREADD.AD<0> ;
  wire \DSP_PREADD.AD<10> ;
  wire \DSP_PREADD.AD<11> ;
  wire \DSP_PREADD.AD<12> ;
  wire \DSP_PREADD.AD<13> ;
  wire \DSP_PREADD.AD<14> ;
  wire \DSP_PREADD.AD<15> ;
  wire \DSP_PREADD.AD<16> ;
  wire \DSP_PREADD.AD<17> ;
  wire \DSP_PREADD.AD<18> ;
  wire \DSP_PREADD.AD<19> ;
  wire \DSP_PREADD.AD<1> ;
  wire \DSP_PREADD.AD<20> ;
  wire \DSP_PREADD.AD<21> ;
  wire \DSP_PREADD.AD<22> ;
  wire \DSP_PREADD.AD<23> ;
  wire \DSP_PREADD.AD<24> ;
  wire \DSP_PREADD.AD<25> ;
  wire \DSP_PREADD.AD<26> ;
  wire \DSP_PREADD.AD<2> ;
  wire \DSP_PREADD.AD<3> ;
  wire \DSP_PREADD.AD<4> ;
  wire \DSP_PREADD.AD<5> ;
  wire \DSP_PREADD.AD<6> ;
  wire \DSP_PREADD.AD<7> ;
  wire \DSP_PREADD.AD<8> ;
  wire \DSP_PREADD.AD<9> ;
  wire \DSP_PREADD_DATA.A2A1<0> ;
  wire \DSP_PREADD_DATA.A2A1<10> ;
  wire \DSP_PREADD_DATA.A2A1<11> ;
  wire \DSP_PREADD_DATA.A2A1<12> ;
  wire \DSP_PREADD_DATA.A2A1<13> ;
  wire \DSP_PREADD_DATA.A2A1<14> ;
  wire \DSP_PREADD_DATA.A2A1<15> ;
  wire \DSP_PREADD_DATA.A2A1<16> ;
  wire \DSP_PREADD_DATA.A2A1<17> ;
  wire \DSP_PREADD_DATA.A2A1<18> ;
  wire \DSP_PREADD_DATA.A2A1<19> ;
  wire \DSP_PREADD_DATA.A2A1<1> ;
  wire \DSP_PREADD_DATA.A2A1<20> ;
  wire \DSP_PREADD_DATA.A2A1<21> ;
  wire \DSP_PREADD_DATA.A2A1<22> ;
  wire \DSP_PREADD_DATA.A2A1<23> ;
  wire \DSP_PREADD_DATA.A2A1<24> ;
  wire \DSP_PREADD_DATA.A2A1<25> ;
  wire \DSP_PREADD_DATA.A2A1<26> ;
  wire \DSP_PREADD_DATA.A2A1<2> ;
  wire \DSP_PREADD_DATA.A2A1<3> ;
  wire \DSP_PREADD_DATA.A2A1<4> ;
  wire \DSP_PREADD_DATA.A2A1<5> ;
  wire \DSP_PREADD_DATA.A2A1<6> ;
  wire \DSP_PREADD_DATA.A2A1<7> ;
  wire \DSP_PREADD_DATA.A2A1<8> ;
  wire \DSP_PREADD_DATA.A2A1<9> ;
  wire \DSP_PREADD_DATA.ADDSUB ;
  wire \DSP_PREADD_DATA.AD_DATA<0> ;
  wire \DSP_PREADD_DATA.AD_DATA<10> ;
  wire \DSP_PREADD_DATA.AD_DATA<11> ;
  wire \DSP_PREADD_DATA.AD_DATA<12> ;
  wire \DSP_PREADD_DATA.AD_DATA<13> ;
  wire \DSP_PREADD_DATA.AD_DATA<14> ;
  wire \DSP_PREADD_DATA.AD_DATA<15> ;
  wire \DSP_PREADD_DATA.AD_DATA<16> ;
  wire \DSP_PREADD_DATA.AD_DATA<17> ;
  wire \DSP_PREADD_DATA.AD_DATA<18> ;
  wire \DSP_PREADD_DATA.AD_DATA<19> ;
  wire \DSP_PREADD_DATA.AD_DATA<1> ;
  wire \DSP_PREADD_DATA.AD_DATA<20> ;
  wire \DSP_PREADD_DATA.AD_DATA<21> ;
  wire \DSP_PREADD_DATA.AD_DATA<22> ;
  wire \DSP_PREADD_DATA.AD_DATA<23> ;
  wire \DSP_PREADD_DATA.AD_DATA<24> ;
  wire \DSP_PREADD_DATA.AD_DATA<25> ;
  wire \DSP_PREADD_DATA.AD_DATA<26> ;
  wire \DSP_PREADD_DATA.AD_DATA<2> ;
  wire \DSP_PREADD_DATA.AD_DATA<3> ;
  wire \DSP_PREADD_DATA.AD_DATA<4> ;
  wire \DSP_PREADD_DATA.AD_DATA<5> ;
  wire \DSP_PREADD_DATA.AD_DATA<6> ;
  wire \DSP_PREADD_DATA.AD_DATA<7> ;
  wire \DSP_PREADD_DATA.AD_DATA<8> ;
  wire \DSP_PREADD_DATA.AD_DATA<9> ;
  wire \DSP_PREADD_DATA.B2B1<0> ;
  wire \DSP_PREADD_DATA.B2B1<10> ;
  wire \DSP_PREADD_DATA.B2B1<11> ;
  wire \DSP_PREADD_DATA.B2B1<12> ;
  wire \DSP_PREADD_DATA.B2B1<13> ;
  wire \DSP_PREADD_DATA.B2B1<14> ;
  wire \DSP_PREADD_DATA.B2B1<15> ;
  wire \DSP_PREADD_DATA.B2B1<16> ;
  wire \DSP_PREADD_DATA.B2B1<17> ;
  wire \DSP_PREADD_DATA.B2B1<1> ;
  wire \DSP_PREADD_DATA.B2B1<2> ;
  wire \DSP_PREADD_DATA.B2B1<3> ;
  wire \DSP_PREADD_DATA.B2B1<4> ;
  wire \DSP_PREADD_DATA.B2B1<5> ;
  wire \DSP_PREADD_DATA.B2B1<6> ;
  wire \DSP_PREADD_DATA.B2B1<7> ;
  wire \DSP_PREADD_DATA.B2B1<8> ;
  wire \DSP_PREADD_DATA.B2B1<9> ;
  wire \DSP_PREADD_DATA.D_DATA<0> ;
  wire \DSP_PREADD_DATA.D_DATA<10> ;
  wire \DSP_PREADD_DATA.D_DATA<11> ;
  wire \DSP_PREADD_DATA.D_DATA<12> ;
  wire \DSP_PREADD_DATA.D_DATA<13> ;
  wire \DSP_PREADD_DATA.D_DATA<14> ;
  wire \DSP_PREADD_DATA.D_DATA<15> ;
  wire \DSP_PREADD_DATA.D_DATA<16> ;
  wire \DSP_PREADD_DATA.D_DATA<17> ;
  wire \DSP_PREADD_DATA.D_DATA<18> ;
  wire \DSP_PREADD_DATA.D_DATA<19> ;
  wire \DSP_PREADD_DATA.D_DATA<1> ;
  wire \DSP_PREADD_DATA.D_DATA<20> ;
  wire \DSP_PREADD_DATA.D_DATA<21> ;
  wire \DSP_PREADD_DATA.D_DATA<22> ;
  wire \DSP_PREADD_DATA.D_DATA<23> ;
  wire \DSP_PREADD_DATA.D_DATA<24> ;
  wire \DSP_PREADD_DATA.D_DATA<25> ;
  wire \DSP_PREADD_DATA.D_DATA<26> ;
  wire \DSP_PREADD_DATA.D_DATA<2> ;
  wire \DSP_PREADD_DATA.D_DATA<3> ;
  wire \DSP_PREADD_DATA.D_DATA<4> ;
  wire \DSP_PREADD_DATA.D_DATA<5> ;
  wire \DSP_PREADD_DATA.D_DATA<6> ;
  wire \DSP_PREADD_DATA.D_DATA<7> ;
  wire \DSP_PREADD_DATA.D_DATA<8> ;
  wire \DSP_PREADD_DATA.D_DATA<9> ;
  wire \DSP_PREADD_DATA.INMODE_2 ;
  wire \DSP_PREADD_DATA.PREADD_AB<0> ;
  wire \DSP_PREADD_DATA.PREADD_AB<10> ;
  wire \DSP_PREADD_DATA.PREADD_AB<11> ;
  wire \DSP_PREADD_DATA.PREADD_AB<12> ;
  wire \DSP_PREADD_DATA.PREADD_AB<13> ;
  wire \DSP_PREADD_DATA.PREADD_AB<14> ;
  wire \DSP_PREADD_DATA.PREADD_AB<15> ;
  wire \DSP_PREADD_DATA.PREADD_AB<16> ;
  wire \DSP_PREADD_DATA.PREADD_AB<17> ;
  wire \DSP_PREADD_DATA.PREADD_AB<18> ;
  wire \DSP_PREADD_DATA.PREADD_AB<19> ;
  wire \DSP_PREADD_DATA.PREADD_AB<1> ;
  wire \DSP_PREADD_DATA.PREADD_AB<20> ;
  wire \DSP_PREADD_DATA.PREADD_AB<21> ;
  wire \DSP_PREADD_DATA.PREADD_AB<22> ;
  wire \DSP_PREADD_DATA.PREADD_AB<23> ;
  wire \DSP_PREADD_DATA.PREADD_AB<24> ;
  wire \DSP_PREADD_DATA.PREADD_AB<25> ;
  wire \DSP_PREADD_DATA.PREADD_AB<26> ;
  wire \DSP_PREADD_DATA.PREADD_AB<2> ;
  wire \DSP_PREADD_DATA.PREADD_AB<3> ;
  wire \DSP_PREADD_DATA.PREADD_AB<4> ;
  wire \DSP_PREADD_DATA.PREADD_AB<5> ;
  wire \DSP_PREADD_DATA.PREADD_AB<6> ;
  wire \DSP_PREADD_DATA.PREADD_AB<7> ;
  wire \DSP_PREADD_DATA.PREADD_AB<8> ;
  wire \DSP_PREADD_DATA.PREADD_AB<9> ;
  wire \D[0] ;
  wire \D[10] ;
  wire \D[11] ;
  wire \D[12] ;
  wire \D[13] ;
  wire \D[14] ;
  wire \D[15] ;
  wire \D[16] ;
  wire \D[17] ;
  wire \D[18] ;
  wire \D[19] ;
  wire \D[1] ;
  wire \D[20] ;
  wire \D[21] ;
  wire \D[22] ;
  wire \D[23] ;
  wire \D[24] ;
  wire \D[25] ;
  wire \D[26] ;
  wire \D[2] ;
  wire \D[3] ;
  wire \D[4] ;
  wire \D[5] ;
  wire \D[6] ;
  wire \D[7] ;
  wire \D[8] ;
  wire \D[9] ;
  wire \INMODE[0] ;
  wire \INMODE[1] ;
  wire \INMODE[2] ;
  wire \INMODE[3] ;
  wire \INMODE[4] ;
  wire MULTSIGNIN;
  wire MULTSIGNOUT;
  wire \OPMODE[0] ;
  wire \OPMODE[1] ;
  wire \OPMODE[2] ;
  wire \OPMODE[3] ;
  wire \OPMODE[4] ;
  wire \OPMODE[5] ;
  wire \OPMODE[6] ;
  wire \OPMODE[7] ;
  wire \OPMODE[8] ;
  wire OVERFLOW;
  wire PATTERNBDETECT;
  wire PATTERNDETECT;
  wire \PCIN[0] ;
  wire \PCIN[10] ;
  wire \PCIN[11] ;
  wire \PCIN[12] ;
  wire \PCIN[13] ;
  wire \PCIN[14] ;
  wire \PCIN[15] ;
  wire \PCIN[16] ;
  wire \PCIN[17] ;
  wire \PCIN[18] ;
  wire \PCIN[19] ;
  wire \PCIN[1] ;
  wire \PCIN[20] ;
  wire \PCIN[21] ;
  wire \PCIN[22] ;
  wire \PCIN[23] ;
  wire \PCIN[24] ;
  wire \PCIN[25] ;
  wire \PCIN[26] ;
  wire \PCIN[27] ;
  wire \PCIN[28] ;
  wire \PCIN[29] ;
  wire \PCIN[2] ;
  wire \PCIN[30] ;
  wire \PCIN[31] ;
  wire \PCIN[32] ;
  wire \PCIN[33] ;
  wire \PCIN[34] ;
  wire \PCIN[35] ;
  wire \PCIN[36] ;
  wire \PCIN[37] ;
  wire \PCIN[38] ;
  wire \PCIN[39] ;
  wire \PCIN[3] ;
  wire \PCIN[40] ;
  wire \PCIN[41] ;
  wire \PCIN[42] ;
  wire \PCIN[43] ;
  wire \PCIN[44] ;
  wire \PCIN[45] ;
  wire \PCIN[46] ;
  wire \PCIN[47] ;
  wire \PCIN[4] ;
  wire \PCIN[5] ;
  wire \PCIN[6] ;
  wire \PCIN[7] ;
  wire \PCIN[8] ;
  wire \PCIN[9] ;
  wire \PCOUT[0] ;
  wire \PCOUT[10] ;
  wire \PCOUT[11] ;
  wire \PCOUT[12] ;
  wire \PCOUT[13] ;
  wire \PCOUT[14] ;
  wire \PCOUT[15] ;
  wire \PCOUT[16] ;
  wire \PCOUT[17] ;
  wire \PCOUT[18] ;
  wire \PCOUT[19] ;
  wire \PCOUT[1] ;
  wire \PCOUT[20] ;
  wire \PCOUT[21] ;
  wire \PCOUT[22] ;
  wire \PCOUT[23] ;
  wire \PCOUT[24] ;
  wire \PCOUT[25] ;
  wire \PCOUT[26] ;
  wire \PCOUT[27] ;
  wire \PCOUT[28] ;
  wire \PCOUT[29] ;
  wire \PCOUT[2] ;
  wire \PCOUT[30] ;
  wire \PCOUT[31] ;
  wire \PCOUT[32] ;
  wire \PCOUT[33] ;
  wire \PCOUT[34] ;
  wire \PCOUT[35] ;
  wire \PCOUT[36] ;
  wire \PCOUT[37] ;
  wire \PCOUT[38] ;
  wire \PCOUT[39] ;
  wire \PCOUT[3] ;
  wire \PCOUT[40] ;
  wire \PCOUT[41] ;
  wire \PCOUT[42] ;
  wire \PCOUT[43] ;
  wire \PCOUT[44] ;
  wire \PCOUT[45] ;
  wire \PCOUT[46] ;
  wire \PCOUT[47] ;
  wire \PCOUT[4] ;
  wire \PCOUT[5] ;
  wire \PCOUT[6] ;
  wire \PCOUT[7] ;
  wire \PCOUT[8] ;
  wire \PCOUT[9] ;
  wire \P[0] ;
  wire \P[10] ;
  wire \P[11] ;
  wire \P[12] ;
  wire \P[13] ;
  wire \P[14] ;
  wire \P[15] ;
  wire \P[16] ;
  wire \P[17] ;
  wire \P[18] ;
  wire \P[19] ;
  wire \P[1] ;
  wire \P[20] ;
  wire \P[21] ;
  wire \P[22] ;
  wire \P[23] ;
  wire \P[24] ;
  wire \P[25] ;
  wire \P[26] ;
  wire \P[27] ;
  wire \P[28] ;
  wire \P[29] ;
  wire \P[2] ;
  wire \P[30] ;
  wire \P[31] ;
  wire \P[32] ;
  wire \P[33] ;
  wire \P[34] ;
  wire \P[35] ;
  wire \P[36] ;
  wire \P[37] ;
  wire \P[38] ;
  wire \P[39] ;
  wire \P[3] ;
  wire \P[40] ;
  wire \P[41] ;
  wire \P[42] ;
  wire \P[43] ;
  wire \P[44] ;
  wire \P[45] ;
  wire \P[46] ;
  wire \P[47] ;
  wire \P[4] ;
  wire \P[5] ;
  wire \P[6] ;
  wire \P[7] ;
  wire \P[8] ;
  wire \P[9] ;
  wire RSTA;
  wire RSTALLCARRYIN;
  wire RSTALUMODE;
  wire RSTB;
  wire RSTC;
  wire RSTCTRL;
  wire RSTD;
  wire RSTINMODE;
  wire RSTM;
  wire RSTP;
  wire UNDERFLOW;
  wire \XOROUT[0] ;
  wire \XOROUT[1] ;
  wire \XOROUT[2] ;
  wire \XOROUT[3] ;
  wire \XOROUT[4] ;
  wire \XOROUT[5] ;
  wire \XOROUT[6] ;
  wire \XOROUT[7] ;

  assign \ACIN[0]  = ACIN[0];
  assign \ACIN[10]  = ACIN[10];
  assign \ACIN[11]  = ACIN[11];
  assign \ACIN[12]  = ACIN[12];
  assign \ACIN[13]  = ACIN[13];
  assign \ACIN[14]  = ACIN[14];
  assign \ACIN[15]  = ACIN[15];
  assign \ACIN[16]  = ACIN[16];
  assign \ACIN[17]  = ACIN[17];
  assign \ACIN[18]  = ACIN[18];
  assign \ACIN[19]  = ACIN[19];
  assign \ACIN[1]  = ACIN[1];
  assign \ACIN[20]  = ACIN[20];
  assign \ACIN[21]  = ACIN[21];
  assign \ACIN[22]  = ACIN[22];
  assign \ACIN[23]  = ACIN[23];
  assign \ACIN[24]  = ACIN[24];
  assign \ACIN[25]  = ACIN[25];
  assign \ACIN[26]  = ACIN[26];
  assign \ACIN[27]  = ACIN[27];
  assign \ACIN[28]  = ACIN[28];
  assign \ACIN[29]  = ACIN[29];
  assign \ACIN[2]  = ACIN[2];
  assign \ACIN[3]  = ACIN[3];
  assign \ACIN[4]  = ACIN[4];
  assign \ACIN[5]  = ACIN[5];
  assign \ACIN[6]  = ACIN[6];
  assign \ACIN[7]  = ACIN[7];
  assign \ACIN[8]  = ACIN[8];
  assign \ACIN[9]  = ACIN[9];
  assign ACOUT[29] = \ACOUT[29] ;
  assign ACOUT[28] = \ACOUT[28] ;
  assign ACOUT[27] = \ACOUT[27] ;
  assign ACOUT[26] = \ACOUT[26] ;
  assign ACOUT[25] = \ACOUT[25] ;
  assign ACOUT[24] = \ACOUT[24] ;
  assign ACOUT[23] = \ACOUT[23] ;
  assign ACOUT[22] = \ACOUT[22] ;
  assign ACOUT[21] = \ACOUT[21] ;
  assign ACOUT[20] = \ACOUT[20] ;
  assign ACOUT[19] = \ACOUT[19] ;
  assign ACOUT[18] = \ACOUT[18] ;
  assign ACOUT[17] = \ACOUT[17] ;
  assign ACOUT[16] = \ACOUT[16] ;
  assign ACOUT[15] = \ACOUT[15] ;
  assign ACOUT[14] = \ACOUT[14] ;
  assign ACOUT[13] = \ACOUT[13] ;
  assign ACOUT[12] = \ACOUT[12] ;
  assign ACOUT[11] = \ACOUT[11] ;
  assign ACOUT[10] = \ACOUT[10] ;
  assign ACOUT[9] = \ACOUT[9] ;
  assign ACOUT[8] = \ACOUT[8] ;
  assign ACOUT[7] = \ACOUT[7] ;
  assign ACOUT[6] = \ACOUT[6] ;
  assign ACOUT[5] = \ACOUT[5] ;
  assign ACOUT[4] = \ACOUT[4] ;
  assign ACOUT[3] = \ACOUT[3] ;
  assign ACOUT[2] = \ACOUT[2] ;
  assign ACOUT[1] = \ACOUT[1] ;
  assign ACOUT[0] = \ACOUT[0] ;
  assign \ALUMODE[0]  = ALUMODE[0];
  assign \ALUMODE[1]  = ALUMODE[1];
  assign \ALUMODE[2]  = ALUMODE[2];
  assign \ALUMODE[3]  = ALUMODE[3];
  assign \A[0]  = A[0];
  assign \A[10]  = A[10];
  assign \A[11]  = A[11];
  assign \A[12]  = A[12];
  assign \A[13]  = A[13];
  assign \A[14]  = A[14];
  assign \A[15]  = A[15];
  assign \A[16]  = A[16];
  assign \A[17]  = A[17];
  assign \A[18]  = A[18];
  assign \A[19]  = A[19];
  assign \A[1]  = A[1];
  assign \A[20]  = A[20];
  assign \A[21]  = A[21];
  assign \A[22]  = A[22];
  assign \A[23]  = A[23];
  assign \A[24]  = A[24];
  assign \A[25]  = A[25];
  assign \A[26]  = A[26];
  assign \A[27]  = A[27];
  assign \A[28]  = A[28];
  assign \A[29]  = A[29];
  assign \A[2]  = A[2];
  assign \A[3]  = A[3];
  assign \A[4]  = A[4];
  assign \A[5]  = A[5];
  assign \A[6]  = A[6];
  assign \A[7]  = A[7];
  assign \A[8]  = A[8];
  assign \A[9]  = A[9];
  assign \BCIN[0]  = BCIN[0];
  assign \BCIN[10]  = BCIN[10];
  assign \BCIN[11]  = BCIN[11];
  assign \BCIN[12]  = BCIN[12];
  assign \BCIN[13]  = BCIN[13];
  assign \BCIN[14]  = BCIN[14];
  assign \BCIN[15]  = BCIN[15];
  assign \BCIN[16]  = BCIN[16];
  assign \BCIN[17]  = BCIN[17];
  assign \BCIN[1]  = BCIN[1];
  assign \BCIN[2]  = BCIN[2];
  assign \BCIN[3]  = BCIN[3];
  assign \BCIN[4]  = BCIN[4];
  assign \BCIN[5]  = BCIN[5];
  assign \BCIN[6]  = BCIN[6];
  assign \BCIN[7]  = BCIN[7];
  assign \BCIN[8]  = BCIN[8];
  assign \BCIN[9]  = BCIN[9];
  assign BCOUT[17] = \BCOUT[17] ;
  assign BCOUT[16] = \BCOUT[16] ;
  assign BCOUT[15] = \BCOUT[15] ;
  assign BCOUT[14] = \BCOUT[14] ;
  assign BCOUT[13] = \BCOUT[13] ;
  assign BCOUT[12] = \BCOUT[12] ;
  assign BCOUT[11] = \BCOUT[11] ;
  assign BCOUT[10] = \BCOUT[10] ;
  assign BCOUT[9] = \BCOUT[9] ;
  assign BCOUT[8] = \BCOUT[8] ;
  assign BCOUT[7] = \BCOUT[7] ;
  assign BCOUT[6] = \BCOUT[6] ;
  assign BCOUT[5] = \BCOUT[5] ;
  assign BCOUT[4] = \BCOUT[4] ;
  assign BCOUT[3] = \BCOUT[3] ;
  assign BCOUT[2] = \BCOUT[2] ;
  assign BCOUT[1] = \BCOUT[1] ;
  assign BCOUT[0] = \BCOUT[0] ;
  assign \B[0]  = B[0];
  assign \B[10]  = B[10];
  assign \B[11]  = B[11];
  assign \B[12]  = B[12];
  assign \B[13]  = B[13];
  assign \B[14]  = B[14];
  assign \B[15]  = B[15];
  assign \B[16]  = B[16];
  assign \B[17]  = B[17];
  assign \B[1]  = B[1];
  assign \B[2]  = B[2];
  assign \B[3]  = B[3];
  assign \B[4]  = B[4];
  assign \B[5]  = B[5];
  assign \B[6]  = B[6];
  assign \B[7]  = B[7];
  assign \B[8]  = B[8];
  assign \B[9]  = B[9];
  assign \CARRYINSEL[0]  = CARRYINSEL[0];
  assign \CARRYINSEL[1]  = CARRYINSEL[1];
  assign \CARRYINSEL[2]  = CARRYINSEL[2];
  assign CARRYOUT[3] = \CARRYOUT[3] ;
  assign CARRYOUT[2] = \CARRYOUT[2] ;
  assign CARRYOUT[1] = \CARRYOUT[1] ;
  assign CARRYOUT[0] = \CARRYOUT[0] ;
  assign \C[0]  = C[0];
  assign \C[10]  = C[10];
  assign \C[11]  = C[11];
  assign \C[12]  = C[12];
  assign \C[13]  = C[13];
  assign \C[14]  = C[14];
  assign \C[15]  = C[15];
  assign \C[16]  = C[16];
  assign \C[17]  = C[17];
  assign \C[18]  = C[18];
  assign \C[19]  = C[19];
  assign \C[1]  = C[1];
  assign \C[20]  = C[20];
  assign \C[21]  = C[21];
  assign \C[22]  = C[22];
  assign \C[23]  = C[23];
  assign \C[24]  = C[24];
  assign \C[25]  = C[25];
  assign \C[26]  = C[26];
  assign \C[27]  = C[27];
  assign \C[28]  = C[28];
  assign \C[29]  = C[29];
  assign \C[2]  = C[2];
  assign \C[30]  = C[30];
  assign \C[31]  = C[31];
  assign \C[32]  = C[32];
  assign \C[33]  = C[33];
  assign \C[34]  = C[34];
  assign \C[35]  = C[35];
  assign \C[36]  = C[36];
  assign \C[37]  = C[37];
  assign \C[38]  = C[38];
  assign \C[39]  = C[39];
  assign \C[3]  = C[3];
  assign \C[40]  = C[40];
  assign \C[41]  = C[41];
  assign \C[42]  = C[42];
  assign \C[43]  = C[43];
  assign \C[44]  = C[44];
  assign \C[45]  = C[45];
  assign \C[46]  = C[46];
  assign \C[47]  = C[47];
  assign \C[4]  = C[4];
  assign \C[5]  = C[5];
  assign \C[6]  = C[6];
  assign \C[7]  = C[7];
  assign \C[8]  = C[8];
  assign \C[9]  = C[9];
  assign \D[0]  = D[0];
  assign \D[10]  = D[10];
  assign \D[11]  = D[11];
  assign \D[12]  = D[12];
  assign \D[13]  = D[13];
  assign \D[14]  = D[14];
  assign \D[15]  = D[15];
  assign \D[16]  = D[16];
  assign \D[17]  = D[17];
  assign \D[18]  = D[18];
  assign \D[19]  = D[19];
  assign \D[1]  = D[1];
  assign \D[20]  = D[20];
  assign \D[21]  = D[21];
  assign \D[22]  = D[22];
  assign \D[23]  = D[23];
  assign \D[24]  = D[24];
  assign \D[25]  = D[25];
  assign \D[26]  = D[26];
  assign \D[2]  = D[2];
  assign \D[3]  = D[3];
  assign \D[4]  = D[4];
  assign \D[5]  = D[5];
  assign \D[6]  = D[6];
  assign \D[7]  = D[7];
  assign \D[8]  = D[8];
  assign \D[9]  = D[9];
  assign \INMODE[0]  = INMODE[0];
  assign \INMODE[1]  = INMODE[1];
  assign \INMODE[2]  = INMODE[2];
  assign \INMODE[3]  = INMODE[3];
  assign \INMODE[4]  = INMODE[4];
  assign \OPMODE[0]  = OPMODE[0];
  assign \OPMODE[1]  = OPMODE[1];
  assign \OPMODE[2]  = OPMODE[2];
  assign \OPMODE[3]  = OPMODE[3];
  assign \OPMODE[4]  = OPMODE[4];
  assign \OPMODE[5]  = OPMODE[5];
  assign \OPMODE[6]  = OPMODE[6];
  assign \OPMODE[7]  = OPMODE[7];
  assign \OPMODE[8]  = OPMODE[8];
  assign P[47] = \P[47] ;
  assign P[46] = \P[46] ;
  assign P[45] = \P[45] ;
  assign P[44] = \P[44] ;
  assign P[43] = \P[43] ;
  assign P[42] = \P[42] ;
  assign P[41] = \P[41] ;
  assign P[40] = \P[40] ;
  assign P[39] = \P[39] ;
  assign P[38] = \P[38] ;
  assign P[37] = \P[37] ;
  assign P[36] = \P[36] ;
  assign P[35] = \P[35] ;
  assign P[34] = \P[34] ;
  assign P[33] = \P[33] ;
  assign P[32] = \P[32] ;
  assign P[31] = \P[31] ;
  assign P[30] = \P[30] ;
  assign P[29] = \P[29] ;
  assign P[28] = \P[28] ;
  assign P[27] = \P[27] ;
  assign P[26] = \P[26] ;
  assign P[25] = \P[25] ;
  assign P[24] = \P[24] ;
  assign P[23] = \P[23] ;
  assign P[22] = \P[22] ;
  assign P[21] = \P[21] ;
  assign P[20] = \P[20] ;
  assign P[19] = \P[19] ;
  assign P[18] = \P[18] ;
  assign P[17] = \P[17] ;
  assign P[16] = \P[16] ;
  assign P[15] = \P[15] ;
  assign P[14] = \P[14] ;
  assign P[13] = \P[13] ;
  assign P[12] = \P[12] ;
  assign P[11] = \P[11] ;
  assign P[10] = \P[10] ;
  assign P[9] = \P[9] ;
  assign P[8] = \P[8] ;
  assign P[7] = \P[7] ;
  assign P[6] = \P[6] ;
  assign P[5] = \P[5] ;
  assign P[4] = \P[4] ;
  assign P[3] = \P[3] ;
  assign P[2] = \P[2] ;
  assign P[1] = \P[1] ;
  assign P[0] = \P[0] ;
  assign \PCIN[0]  = PCIN[0];
  assign \PCIN[10]  = PCIN[10];
  assign \PCIN[11]  = PCIN[11];
  assign \PCIN[12]  = PCIN[12];
  assign \PCIN[13]  = PCIN[13];
  assign \PCIN[14]  = PCIN[14];
  assign \PCIN[15]  = PCIN[15];
  assign \PCIN[16]  = PCIN[16];
  assign \PCIN[17]  = PCIN[17];
  assign \PCIN[18]  = PCIN[18];
  assign \PCIN[19]  = PCIN[19];
  assign \PCIN[1]  = PCIN[1];
  assign \PCIN[20]  = PCIN[20];
  assign \PCIN[21]  = PCIN[21];
  assign \PCIN[22]  = PCIN[22];
  assign \PCIN[23]  = PCIN[23];
  assign \PCIN[24]  = PCIN[24];
  assign \PCIN[25]  = PCIN[25];
  assign \PCIN[26]  = PCIN[26];
  assign \PCIN[27]  = PCIN[27];
  assign \PCIN[28]  = PCIN[28];
  assign \PCIN[29]  = PCIN[29];
  assign \PCIN[2]  = PCIN[2];
  assign \PCIN[30]  = PCIN[30];
  assign \PCIN[31]  = PCIN[31];
  assign \PCIN[32]  = PCIN[32];
  assign \PCIN[33]  = PCIN[33];
  assign \PCIN[34]  = PCIN[34];
  assign \PCIN[35]  = PCIN[35];
  assign \PCIN[36]  = PCIN[36];
  assign \PCIN[37]  = PCIN[37];
  assign \PCIN[38]  = PCIN[38];
  assign \PCIN[39]  = PCIN[39];
  assign \PCIN[3]  = PCIN[3];
  assign \PCIN[40]  = PCIN[40];
  assign \PCIN[41]  = PCIN[41];
  assign \PCIN[42]  = PCIN[42];
  assign \PCIN[43]  = PCIN[43];
  assign \PCIN[44]  = PCIN[44];
  assign \PCIN[45]  = PCIN[45];
  assign \PCIN[46]  = PCIN[46];
  assign \PCIN[47]  = PCIN[47];
  assign \PCIN[4]  = PCIN[4];
  assign \PCIN[5]  = PCIN[5];
  assign \PCIN[6]  = PCIN[6];
  assign \PCIN[7]  = PCIN[7];
  assign \PCIN[8]  = PCIN[8];
  assign \PCIN[9]  = PCIN[9];
  assign PCOUT[47] = \PCOUT[47] ;
  assign PCOUT[46] = \PCOUT[46] ;
  assign PCOUT[45] = \PCOUT[45] ;
  assign PCOUT[44] = \PCOUT[44] ;
  assign PCOUT[43] = \PCOUT[43] ;
  assign PCOUT[42] = \PCOUT[42] ;
  assign PCOUT[41] = \PCOUT[41] ;
  assign PCOUT[40] = \PCOUT[40] ;
  assign PCOUT[39] = \PCOUT[39] ;
  assign PCOUT[38] = \PCOUT[38] ;
  assign PCOUT[37] = \PCOUT[37] ;
  assign PCOUT[36] = \PCOUT[36] ;
  assign PCOUT[35] = \PCOUT[35] ;
  assign PCOUT[34] = \PCOUT[34] ;
  assign PCOUT[33] = \PCOUT[33] ;
  assign PCOUT[32] = \PCOUT[32] ;
  assign PCOUT[31] = \PCOUT[31] ;
  assign PCOUT[30] = \PCOUT[30] ;
  assign PCOUT[29] = \PCOUT[29] ;
  assign PCOUT[28] = \PCOUT[28] ;
  assign PCOUT[27] = \PCOUT[27] ;
  assign PCOUT[26] = \PCOUT[26] ;
  assign PCOUT[25] = \PCOUT[25] ;
  assign PCOUT[24] = \PCOUT[24] ;
  assign PCOUT[23] = \PCOUT[23] ;
  assign PCOUT[22] = \PCOUT[22] ;
  assign PCOUT[21] = \PCOUT[21] ;
  assign PCOUT[20] = \PCOUT[20] ;
  assign PCOUT[19] = \PCOUT[19] ;
  assign PCOUT[18] = \PCOUT[18] ;
  assign PCOUT[17] = \PCOUT[17] ;
  assign PCOUT[16] = \PCOUT[16] ;
  assign PCOUT[15] = \PCOUT[15] ;
  assign PCOUT[14] = \PCOUT[14] ;
  assign PCOUT[13] = \PCOUT[13] ;
  assign PCOUT[12] = \PCOUT[12] ;
  assign PCOUT[11] = \PCOUT[11] ;
  assign PCOUT[10] = \PCOUT[10] ;
  assign PCOUT[9] = \PCOUT[9] ;
  assign PCOUT[8] = \PCOUT[8] ;
  assign PCOUT[7] = \PCOUT[7] ;
  assign PCOUT[6] = \PCOUT[6] ;
  assign PCOUT[5] = \PCOUT[5] ;
  assign PCOUT[4] = \PCOUT[4] ;
  assign PCOUT[3] = \PCOUT[3] ;
  assign PCOUT[2] = \PCOUT[2] ;
  assign PCOUT[1] = \PCOUT[1] ;
  assign PCOUT[0] = \PCOUT[0] ;
  assign XOROUT[7] = \XOROUT[7] ;
  assign XOROUT[6] = \XOROUT[6] ;
  assign XOROUT[5] = \XOROUT[5] ;
  assign XOROUT[4] = \XOROUT[4] ;
  assign XOROUT[3] = \XOROUT[3] ;
  assign XOROUT[2] = \XOROUT[2] ;
  assign XOROUT[1] = \XOROUT[1] ;
  assign XOROUT[0] = \XOROUT[0] ;
  DSP_ALU #(
    .ALUMODEREG(0),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_OPMODE_INVERTED(9'b000000000),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .MREG(0),
    .OPMODEREG(0),
    .RND(48'h000000000000),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")) 
    DSP_ALU_INST
       (.ALUMODE({\ALUMODE[3] ,\ALUMODE[2] ,\ALUMODE[1] ,\ALUMODE[0] }),
        .ALUMODE10(\DSP_ALU.ALUMODE10 ),
        .ALU_OUT({\DSP_ALU.ALU_OUT<47> ,\DSP_ALU.ALU_OUT<46> ,\DSP_ALU.ALU_OUT<45> ,\DSP_ALU.ALU_OUT<44> ,\DSP_ALU.ALU_OUT<43> ,\DSP_ALU.ALU_OUT<42> ,\DSP_ALU.ALU_OUT<41> ,\DSP_ALU.ALU_OUT<40> ,\DSP_ALU.ALU_OUT<39> ,\DSP_ALU.ALU_OUT<38> ,\DSP_ALU.ALU_OUT<37> ,\DSP_ALU.ALU_OUT<36> ,\DSP_ALU.ALU_OUT<35> ,\DSP_ALU.ALU_OUT<34> ,\DSP_ALU.ALU_OUT<33> ,\DSP_ALU.ALU_OUT<32> ,\DSP_ALU.ALU_OUT<31> ,\DSP_ALU.ALU_OUT<30> ,\DSP_ALU.ALU_OUT<29> ,\DSP_ALU.ALU_OUT<28> ,\DSP_ALU.ALU_OUT<27> ,\DSP_ALU.ALU_OUT<26> ,\DSP_ALU.ALU_OUT<25> ,\DSP_ALU.ALU_OUT<24> ,\DSP_ALU.ALU_OUT<23> ,\DSP_ALU.ALU_OUT<22> ,\DSP_ALU.ALU_OUT<21> ,\DSP_ALU.ALU_OUT<20> ,\DSP_ALU.ALU_OUT<19> ,\DSP_ALU.ALU_OUT<18> ,\DSP_ALU.ALU_OUT<17> ,\DSP_ALU.ALU_OUT<16> ,\DSP_ALU.ALU_OUT<15> ,\DSP_ALU.ALU_OUT<14> ,\DSP_ALU.ALU_OUT<13> ,\DSP_ALU.ALU_OUT<12> ,\DSP_ALU.ALU_OUT<11> ,\DSP_ALU.ALU_OUT<10> ,\DSP_ALU.ALU_OUT<9> ,\DSP_ALU.ALU_OUT<8> ,\DSP_ALU.ALU_OUT<7> ,\DSP_ALU.ALU_OUT<6> ,\DSP_ALU.ALU_OUT<5> ,\DSP_ALU.ALU_OUT<4> ,\DSP_ALU.ALU_OUT<3> ,\DSP_ALU.ALU_OUT<2> ,\DSP_ALU.ALU_OUT<1> ,\DSP_ALU.ALU_OUT<0> }),
        .AMULT26(\DSP_MULTIPLIER.AMULT26 ),
        .A_ALU({\DSP_A_B_DATA.A_ALU<29> ,\DSP_A_B_DATA.A_ALU<28> ,\DSP_A_B_DATA.A_ALU<27> ,\DSP_A_B_DATA.A_ALU<26> ,\DSP_A_B_DATA.A_ALU<25> ,\DSP_A_B_DATA.A_ALU<24> ,\DSP_A_B_DATA.A_ALU<23> ,\DSP_A_B_DATA.A_ALU<22> ,\DSP_A_B_DATA.A_ALU<21> ,\DSP_A_B_DATA.A_ALU<20> ,\DSP_A_B_DATA.A_ALU<19> ,\DSP_A_B_DATA.A_ALU<18> ,\DSP_A_B_DATA.A_ALU<17> ,\DSP_A_B_DATA.A_ALU<16> ,\DSP_A_B_DATA.A_ALU<15> ,\DSP_A_B_DATA.A_ALU<14> ,\DSP_A_B_DATA.A_ALU<13> ,\DSP_A_B_DATA.A_ALU<12> ,\DSP_A_B_DATA.A_ALU<11> ,\DSP_A_B_DATA.A_ALU<10> ,\DSP_A_B_DATA.A_ALU<9> ,\DSP_A_B_DATA.A_ALU<8> ,\DSP_A_B_DATA.A_ALU<7> ,\DSP_A_B_DATA.A_ALU<6> ,\DSP_A_B_DATA.A_ALU<5> ,\DSP_A_B_DATA.A_ALU<4> ,\DSP_A_B_DATA.A_ALU<3> ,\DSP_A_B_DATA.A_ALU<2> ,\DSP_A_B_DATA.A_ALU<1> ,\DSP_A_B_DATA.A_ALU<0> }),
        .BMULT17(\DSP_MULTIPLIER.BMULT17 ),
        .B_ALU({\DSP_A_B_DATA.B_ALU<17> ,\DSP_A_B_DATA.B_ALU<16> ,\DSP_A_B_DATA.B_ALU<15> ,\DSP_A_B_DATA.B_ALU<14> ,\DSP_A_B_DATA.B_ALU<13> ,\DSP_A_B_DATA.B_ALU<12> ,\DSP_A_B_DATA.B_ALU<11> ,\DSP_A_B_DATA.B_ALU<10> ,\DSP_A_B_DATA.B_ALU<9> ,\DSP_A_B_DATA.B_ALU<8> ,\DSP_A_B_DATA.B_ALU<7> ,\DSP_A_B_DATA.B_ALU<6> ,\DSP_A_B_DATA.B_ALU<5> ,\DSP_A_B_DATA.B_ALU<4> ,\DSP_A_B_DATA.B_ALU<3> ,\DSP_A_B_DATA.B_ALU<2> ,\DSP_A_B_DATA.B_ALU<1> ,\DSP_A_B_DATA.B_ALU<0> }),
        .CARRYCASCIN(CARRYCASCIN),
        .CARRYIN(CARRYIN),
        .CARRYINSEL({\CARRYINSEL[2] ,\CARRYINSEL[1] ,\CARRYINSEL[0] }),
        .CCOUT(\DSP_OUTPUT.CCOUT_FB ),
        .CEALUMODE(CEALUMODE),
        .CECARRYIN(CECARRYIN),
        .CECTRL(CECTRL),
        .CEM(CEM),
        .CLK(CLK),
        .COUT({\DSP_ALU.COUT<3> ,\DSP_ALU.COUT<2> ,\DSP_ALU.COUT<1> ,\DSP_ALU.COUT<0> }),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .MULTSIGNIN(MULTSIGNIN),
        .MULTSIGN_ALU(\DSP_ALU.MULTSIGN_ALU ),
        .OPMODE({\OPMODE[8] ,\OPMODE[7] ,\OPMODE[6] ,\OPMODE[5] ,\OPMODE[4] ,\OPMODE[3] ,\OPMODE[2] ,\OPMODE[1] ,\OPMODE[0] }),
        .PCIN({\PCIN[47] ,\PCIN[46] ,\PCIN[45] ,\PCIN[44] ,\PCIN[43] ,\PCIN[42] ,\PCIN[41] ,\PCIN[40] ,\PCIN[39] ,\PCIN[38] ,\PCIN[37] ,\PCIN[36] ,\PCIN[35] ,\PCIN[34] ,\PCIN[33] ,\PCIN[32] ,\PCIN[31] ,\PCIN[30] ,\PCIN[29] ,\PCIN[28] ,\PCIN[27] ,\PCIN[26] ,\PCIN[25] ,\PCIN[24] ,\PCIN[23] ,\PCIN[22] ,\PCIN[21] ,\PCIN[20] ,\PCIN[19] ,\PCIN[18] ,\PCIN[17] ,\PCIN[16] ,\PCIN[15] ,\PCIN[14] ,\PCIN[13] ,\PCIN[12] ,\PCIN[11] ,\PCIN[10] ,\PCIN[9] ,\PCIN[8] ,\PCIN[7] ,\PCIN[6] ,\PCIN[5] ,\PCIN[4] ,\PCIN[3] ,\PCIN[2] ,\PCIN[1] ,\PCIN[0] }),
        .P_FDBK({\DSP_OUTPUT.P_FDBK<47> ,\DSP_OUTPUT.P_FDBK<46> ,\DSP_OUTPUT.P_FDBK<45> ,\DSP_OUTPUT.P_FDBK<44> ,\DSP_OUTPUT.P_FDBK<43> ,\DSP_OUTPUT.P_FDBK<42> ,\DSP_OUTPUT.P_FDBK<41> ,\DSP_OUTPUT.P_FDBK<40> ,\DSP_OUTPUT.P_FDBK<39> ,\DSP_OUTPUT.P_FDBK<38> ,\DSP_OUTPUT.P_FDBK<37> ,\DSP_OUTPUT.P_FDBK<36> ,\DSP_OUTPUT.P_FDBK<35> ,\DSP_OUTPUT.P_FDBK<34> ,\DSP_OUTPUT.P_FDBK<33> ,\DSP_OUTPUT.P_FDBK<32> ,\DSP_OUTPUT.P_FDBK<31> ,\DSP_OUTPUT.P_FDBK<30> ,\DSP_OUTPUT.P_FDBK<29> ,\DSP_OUTPUT.P_FDBK<28> ,\DSP_OUTPUT.P_FDBK<27> ,\DSP_OUTPUT.P_FDBK<26> ,\DSP_OUTPUT.P_FDBK<25> ,\DSP_OUTPUT.P_FDBK<24> ,\DSP_OUTPUT.P_FDBK<23> ,\DSP_OUTPUT.P_FDBK<22> ,\DSP_OUTPUT.P_FDBK<21> ,\DSP_OUTPUT.P_FDBK<20> ,\DSP_OUTPUT.P_FDBK<19> ,\DSP_OUTPUT.P_FDBK<18> ,\DSP_OUTPUT.P_FDBK<17> ,\DSP_OUTPUT.P_FDBK<16> ,\DSP_OUTPUT.P_FDBK<15> ,\DSP_OUTPUT.P_FDBK<14> ,\DSP_OUTPUT.P_FDBK<13> ,\DSP_OUTPUT.P_FDBK<12> ,\DSP_OUTPUT.P_FDBK<11> ,\DSP_OUTPUT.P_FDBK<10> ,\DSP_OUTPUT.P_FDBK<9> ,\DSP_OUTPUT.P_FDBK<8> ,\DSP_OUTPUT.P_FDBK<7> ,\DSP_OUTPUT.P_FDBK<6> ,\DSP_OUTPUT.P_FDBK<5> ,\DSP_OUTPUT.P_FDBK<4> ,\DSP_OUTPUT.P_FDBK<3> ,\DSP_OUTPUT.P_FDBK<2> ,\DSP_OUTPUT.P_FDBK<1> ,\DSP_OUTPUT.P_FDBK<0> }),
        .P_FDBK_47(\DSP_OUTPUT.P_FDBK_47 ),
        .RSTALLCARRYIN(RSTALLCARRYIN),
        .RSTALUMODE(RSTALUMODE),
        .RSTCTRL(RSTCTRL),
        .U_DATA({\DSP_M_DATA.U_DATA<44> ,\DSP_M_DATA.U_DATA<43> ,\DSP_M_DATA.U_DATA<42> ,\DSP_M_DATA.U_DATA<41> ,\DSP_M_DATA.U_DATA<40> ,\DSP_M_DATA.U_DATA<39> ,\DSP_M_DATA.U_DATA<38> ,\DSP_M_DATA.U_DATA<37> ,\DSP_M_DATA.U_DATA<36> ,\DSP_M_DATA.U_DATA<35> ,\DSP_M_DATA.U_DATA<34> ,\DSP_M_DATA.U_DATA<33> ,\DSP_M_DATA.U_DATA<32> ,\DSP_M_DATA.U_DATA<31> ,\DSP_M_DATA.U_DATA<30> ,\DSP_M_DATA.U_DATA<29> ,\DSP_M_DATA.U_DATA<28> ,\DSP_M_DATA.U_DATA<27> ,\DSP_M_DATA.U_DATA<26> ,\DSP_M_DATA.U_DATA<25> ,\DSP_M_DATA.U_DATA<24> ,\DSP_M_DATA.U_DATA<23> ,\DSP_M_DATA.U_DATA<22> ,\DSP_M_DATA.U_DATA<21> ,\DSP_M_DATA.U_DATA<20> ,\DSP_M_DATA.U_DATA<19> ,\DSP_M_DATA.U_DATA<18> ,\DSP_M_DATA.U_DATA<17> ,\DSP_M_DATA.U_DATA<16> ,\DSP_M_DATA.U_DATA<15> ,\DSP_M_DATA.U_DATA<14> ,\DSP_M_DATA.U_DATA<13> ,\DSP_M_DATA.U_DATA<12> ,\DSP_M_DATA.U_DATA<11> ,\DSP_M_DATA.U_DATA<10> ,\DSP_M_DATA.U_DATA<9> ,\DSP_M_DATA.U_DATA<8> ,\DSP_M_DATA.U_DATA<7> ,\DSP_M_DATA.U_DATA<6> ,\DSP_M_DATA.U_DATA<5> ,\DSP_M_DATA.U_DATA<4> ,\DSP_M_DATA.U_DATA<3> ,\DSP_M_DATA.U_DATA<2> ,\DSP_M_DATA.U_DATA<1> ,\DSP_M_DATA.U_DATA<0> }),
        .V_DATA({\DSP_M_DATA.V_DATA<44> ,\DSP_M_DATA.V_DATA<43> ,\DSP_M_DATA.V_DATA<42> ,\DSP_M_DATA.V_DATA<41> ,\DSP_M_DATA.V_DATA<40> ,\DSP_M_DATA.V_DATA<39> ,\DSP_M_DATA.V_DATA<38> ,\DSP_M_DATA.V_DATA<37> ,\DSP_M_DATA.V_DATA<36> ,\DSP_M_DATA.V_DATA<35> ,\DSP_M_DATA.V_DATA<34> ,\DSP_M_DATA.V_DATA<33> ,\DSP_M_DATA.V_DATA<32> ,\DSP_M_DATA.V_DATA<31> ,\DSP_M_DATA.V_DATA<30> ,\DSP_M_DATA.V_DATA<29> ,\DSP_M_DATA.V_DATA<28> ,\DSP_M_DATA.V_DATA<27> ,\DSP_M_DATA.V_DATA<26> ,\DSP_M_DATA.V_DATA<25> ,\DSP_M_DATA.V_DATA<24> ,\DSP_M_DATA.V_DATA<23> ,\DSP_M_DATA.V_DATA<22> ,\DSP_M_DATA.V_DATA<21> ,\DSP_M_DATA.V_DATA<20> ,\DSP_M_DATA.V_DATA<19> ,\DSP_M_DATA.V_DATA<18> ,\DSP_M_DATA.V_DATA<17> ,\DSP_M_DATA.V_DATA<16> ,\DSP_M_DATA.V_DATA<15> ,\DSP_M_DATA.V_DATA<14> ,\DSP_M_DATA.V_DATA<13> ,\DSP_M_DATA.V_DATA<12> ,\DSP_M_DATA.V_DATA<11> ,\DSP_M_DATA.V_DATA<10> ,\DSP_M_DATA.V_DATA<9> ,\DSP_M_DATA.V_DATA<8> ,\DSP_M_DATA.V_DATA<7> ,\DSP_M_DATA.V_DATA<6> ,\DSP_M_DATA.V_DATA<5> ,\DSP_M_DATA.V_DATA<4> ,\DSP_M_DATA.V_DATA<3> ,\DSP_M_DATA.V_DATA<2> ,\DSP_M_DATA.V_DATA<1> ,\DSP_M_DATA.V_DATA<0> }),
        .XOR_MX({\DSP_ALU.XOR_MX<7> ,\DSP_ALU.XOR_MX<6> ,\DSP_ALU.XOR_MX<5> ,\DSP_ALU.XOR_MX<4> ,\DSP_ALU.XOR_MX<3> ,\DSP_ALU.XOR_MX<2> ,\DSP_ALU.XOR_MX<1> ,\DSP_ALU.XOR_MX<0> }));
  DSP_A_B_DATA #(
    .ACASCREG(0),
    .AREG(0),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0)) 
    DSP_A_B_DATA_INST
       (.A({\A[29] ,\A[28] ,\A[27] ,\A[26] ,\A[25] ,\A[24] ,\A[23] ,\A[22] ,\A[21] ,\A[20] ,\A[19] ,\A[18] ,\A[17] ,\A[16] ,\A[15] ,\A[14] ,\A[13] ,\A[12] ,\A[11] ,\A[10] ,\A[9] ,\A[8] ,\A[7] ,\A[6] ,\A[5] ,\A[4] ,\A[3] ,\A[2] ,\A[1] ,\A[0] }),
        .A1_DATA({\DSP_A_B_DATA.A1_DATA<26> ,\DSP_A_B_DATA.A1_DATA<25> ,\DSP_A_B_DATA.A1_DATA<24> ,\DSP_A_B_DATA.A1_DATA<23> ,\DSP_A_B_DATA.A1_DATA<22> ,\DSP_A_B_DATA.A1_DATA<21> ,\DSP_A_B_DATA.A1_DATA<20> ,\DSP_A_B_DATA.A1_DATA<19> ,\DSP_A_B_DATA.A1_DATA<18> ,\DSP_A_B_DATA.A1_DATA<17> ,\DSP_A_B_DATA.A1_DATA<16> ,\DSP_A_B_DATA.A1_DATA<15> ,\DSP_A_B_DATA.A1_DATA<14> ,\DSP_A_B_DATA.A1_DATA<13> ,\DSP_A_B_DATA.A1_DATA<12> ,\DSP_A_B_DATA.A1_DATA<11> ,\DSP_A_B_DATA.A1_DATA<10> ,\DSP_A_B_DATA.A1_DATA<9> ,\DSP_A_B_DATA.A1_DATA<8> ,\DSP_A_B_DATA.A1_DATA<7> ,\DSP_A_B_DATA.A1_DATA<6> ,\DSP_A_B_DATA.A1_DATA<5> ,\DSP_A_B_DATA.A1_DATA<4> ,\DSP_A_B_DATA.A1_DATA<3> ,\DSP_A_B_DATA.A1_DATA<2> ,\DSP_A_B_DATA.A1_DATA<1> ,\DSP_A_B_DATA.A1_DATA<0> }),
        .A2_DATA({\DSP_A_B_DATA.A2_DATA<26> ,\DSP_A_B_DATA.A2_DATA<25> ,\DSP_A_B_DATA.A2_DATA<24> ,\DSP_A_B_DATA.A2_DATA<23> ,\DSP_A_B_DATA.A2_DATA<22> ,\DSP_A_B_DATA.A2_DATA<21> ,\DSP_A_B_DATA.A2_DATA<20> ,\DSP_A_B_DATA.A2_DATA<19> ,\DSP_A_B_DATA.A2_DATA<18> ,\DSP_A_B_DATA.A2_DATA<17> ,\DSP_A_B_DATA.A2_DATA<16> ,\DSP_A_B_DATA.A2_DATA<15> ,\DSP_A_B_DATA.A2_DATA<14> ,\DSP_A_B_DATA.A2_DATA<13> ,\DSP_A_B_DATA.A2_DATA<12> ,\DSP_A_B_DATA.A2_DATA<11> ,\DSP_A_B_DATA.A2_DATA<10> ,\DSP_A_B_DATA.A2_DATA<9> ,\DSP_A_B_DATA.A2_DATA<8> ,\DSP_A_B_DATA.A2_DATA<7> ,\DSP_A_B_DATA.A2_DATA<6> ,\DSP_A_B_DATA.A2_DATA<5> ,\DSP_A_B_DATA.A2_DATA<4> ,\DSP_A_B_DATA.A2_DATA<3> ,\DSP_A_B_DATA.A2_DATA<2> ,\DSP_A_B_DATA.A2_DATA<1> ,\DSP_A_B_DATA.A2_DATA<0> }),
        .ACIN({\ACIN[29] ,\ACIN[28] ,\ACIN[27] ,\ACIN[26] ,\ACIN[25] ,\ACIN[24] ,\ACIN[23] ,\ACIN[22] ,\ACIN[21] ,\ACIN[20] ,\ACIN[19] ,\ACIN[18] ,\ACIN[17] ,\ACIN[16] ,\ACIN[15] ,\ACIN[14] ,\ACIN[13] ,\ACIN[12] ,\ACIN[11] ,\ACIN[10] ,\ACIN[9] ,\ACIN[8] ,\ACIN[7] ,\ACIN[6] ,\ACIN[5] ,\ACIN[4] ,\ACIN[3] ,\ACIN[2] ,\ACIN[1] ,\ACIN[0] }),
        .ACOUT({\ACOUT[29] ,\ACOUT[28] ,\ACOUT[27] ,\ACOUT[26] ,\ACOUT[25] ,\ACOUT[24] ,\ACOUT[23] ,\ACOUT[22] ,\ACOUT[21] ,\ACOUT[20] ,\ACOUT[19] ,\ACOUT[18] ,\ACOUT[17] ,\ACOUT[16] ,\ACOUT[15] ,\ACOUT[14] ,\ACOUT[13] ,\ACOUT[12] ,\ACOUT[11] ,\ACOUT[10] ,\ACOUT[9] ,\ACOUT[8] ,\ACOUT[7] ,\ACOUT[6] ,\ACOUT[5] ,\ACOUT[4] ,\ACOUT[3] ,\ACOUT[2] ,\ACOUT[1] ,\ACOUT[0] }),
        .A_ALU({\DSP_A_B_DATA.A_ALU<29> ,\DSP_A_B_DATA.A_ALU<28> ,\DSP_A_B_DATA.A_ALU<27> ,\DSP_A_B_DATA.A_ALU<26> ,\DSP_A_B_DATA.A_ALU<25> ,\DSP_A_B_DATA.A_ALU<24> ,\DSP_A_B_DATA.A_ALU<23> ,\DSP_A_B_DATA.A_ALU<22> ,\DSP_A_B_DATA.A_ALU<21> ,\DSP_A_B_DATA.A_ALU<20> ,\DSP_A_B_DATA.A_ALU<19> ,\DSP_A_B_DATA.A_ALU<18> ,\DSP_A_B_DATA.A_ALU<17> ,\DSP_A_B_DATA.A_ALU<16> ,\DSP_A_B_DATA.A_ALU<15> ,\DSP_A_B_DATA.A_ALU<14> ,\DSP_A_B_DATA.A_ALU<13> ,\DSP_A_B_DATA.A_ALU<12> ,\DSP_A_B_DATA.A_ALU<11> ,\DSP_A_B_DATA.A_ALU<10> ,\DSP_A_B_DATA.A_ALU<9> ,\DSP_A_B_DATA.A_ALU<8> ,\DSP_A_B_DATA.A_ALU<7> ,\DSP_A_B_DATA.A_ALU<6> ,\DSP_A_B_DATA.A_ALU<5> ,\DSP_A_B_DATA.A_ALU<4> ,\DSP_A_B_DATA.A_ALU<3> ,\DSP_A_B_DATA.A_ALU<2> ,\DSP_A_B_DATA.A_ALU<1> ,\DSP_A_B_DATA.A_ALU<0> }),
        .B({\B[17] ,\B[16] ,\B[15] ,\B[14] ,\B[13] ,\B[12] ,\B[11] ,\B[10] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,\B[0] }),
        .B1_DATA({\DSP_A_B_DATA.B1_DATA<17> ,\DSP_A_B_DATA.B1_DATA<16> ,\DSP_A_B_DATA.B1_DATA<15> ,\DSP_A_B_DATA.B1_DATA<14> ,\DSP_A_B_DATA.B1_DATA<13> ,\DSP_A_B_DATA.B1_DATA<12> ,\DSP_A_B_DATA.B1_DATA<11> ,\DSP_A_B_DATA.B1_DATA<10> ,\DSP_A_B_DATA.B1_DATA<9> ,\DSP_A_B_DATA.B1_DATA<8> ,\DSP_A_B_DATA.B1_DATA<7> ,\DSP_A_B_DATA.B1_DATA<6> ,\DSP_A_B_DATA.B1_DATA<5> ,\DSP_A_B_DATA.B1_DATA<4> ,\DSP_A_B_DATA.B1_DATA<3> ,\DSP_A_B_DATA.B1_DATA<2> ,\DSP_A_B_DATA.B1_DATA<1> ,\DSP_A_B_DATA.B1_DATA<0> }),
        .B2_DATA({\DSP_A_B_DATA.B2_DATA<17> ,\DSP_A_B_DATA.B2_DATA<16> ,\DSP_A_B_DATA.B2_DATA<15> ,\DSP_A_B_DATA.B2_DATA<14> ,\DSP_A_B_DATA.B2_DATA<13> ,\DSP_A_B_DATA.B2_DATA<12> ,\DSP_A_B_DATA.B2_DATA<11> ,\DSP_A_B_DATA.B2_DATA<10> ,\DSP_A_B_DATA.B2_DATA<9> ,\DSP_A_B_DATA.B2_DATA<8> ,\DSP_A_B_DATA.B2_DATA<7> ,\DSP_A_B_DATA.B2_DATA<6> ,\DSP_A_B_DATA.B2_DATA<5> ,\DSP_A_B_DATA.B2_DATA<4> ,\DSP_A_B_DATA.B2_DATA<3> ,\DSP_A_B_DATA.B2_DATA<2> ,\DSP_A_B_DATA.B2_DATA<1> ,\DSP_A_B_DATA.B2_DATA<0> }),
        .BCIN({\BCIN[17] ,\BCIN[16] ,\BCIN[15] ,\BCIN[14] ,\BCIN[13] ,\BCIN[12] ,\BCIN[11] ,\BCIN[10] ,\BCIN[9] ,\BCIN[8] ,\BCIN[7] ,\BCIN[6] ,\BCIN[5] ,\BCIN[4] ,\BCIN[3] ,\BCIN[2] ,\BCIN[1] ,\BCIN[0] }),
        .BCOUT({\BCOUT[17] ,\BCOUT[16] ,\BCOUT[15] ,\BCOUT[14] ,\BCOUT[13] ,\BCOUT[12] ,\BCOUT[11] ,\BCOUT[10] ,\BCOUT[9] ,\BCOUT[8] ,\BCOUT[7] ,\BCOUT[6] ,\BCOUT[5] ,\BCOUT[4] ,\BCOUT[3] ,\BCOUT[2] ,\BCOUT[1] ,\BCOUT[0] }),
        .B_ALU({\DSP_A_B_DATA.B_ALU<17> ,\DSP_A_B_DATA.B_ALU<16> ,\DSP_A_B_DATA.B_ALU<15> ,\DSP_A_B_DATA.B_ALU<14> ,\DSP_A_B_DATA.B_ALU<13> ,\DSP_A_B_DATA.B_ALU<12> ,\DSP_A_B_DATA.B_ALU<11> ,\DSP_A_B_DATA.B_ALU<10> ,\DSP_A_B_DATA.B_ALU<9> ,\DSP_A_B_DATA.B_ALU<8> ,\DSP_A_B_DATA.B_ALU<7> ,\DSP_A_B_DATA.B_ALU<6> ,\DSP_A_B_DATA.B_ALU<5> ,\DSP_A_B_DATA.B_ALU<4> ,\DSP_A_B_DATA.B_ALU<3> ,\DSP_A_B_DATA.B_ALU<2> ,\DSP_A_B_DATA.B_ALU<1> ,\DSP_A_B_DATA.B_ALU<0> }),
        .CEA1(CEA1),
        .CEA2(CEA2),
        .CEB1(CEB1),
        .CEB2(CEB2),
        .CLK(CLK),
        .RSTA(RSTA),
        .RSTB(RSTB));
  DSP_C_DATA #(
    .CREG(0),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0)) 
    DSP_C_DATA_INST
       (.C({\C[47] ,\C[46] ,\C[45] ,\C[44] ,\C[43] ,\C[42] ,\C[41] ,\C[40] ,\C[39] ,\C[38] ,\C[37] ,\C[36] ,\C[35] ,\C[34] ,\C[33] ,\C[32] ,\C[31] ,\C[30] ,\C[29] ,\C[28] ,\C[27] ,\C[26] ,\C[25] ,\C[24] ,\C[23] ,\C[22] ,\C[21] ,\C[20] ,\C[19] ,\C[18] ,\C[17] ,\C[16] ,\C[15] ,\C[14] ,\C[13] ,\C[12] ,\C[11] ,\C[10] ,\C[9] ,\C[8] ,\C[7] ,\C[6] ,\C[5] ,\C[4] ,\C[3] ,\C[2] ,\C[1] ,\C[0] }),
        .CEC(CEC),
        .CLK(CLK),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .RSTC(RSTC));
  DSP_MULTIPLIER #(
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .USE_MULT("MULTIPLY")) 
    DSP_MULTIPLIER_INST
       (.A2A1({\DSP_PREADD_DATA.A2A1<26> ,\DSP_PREADD_DATA.A2A1<25> ,\DSP_PREADD_DATA.A2A1<24> ,\DSP_PREADD_DATA.A2A1<23> ,\DSP_PREADD_DATA.A2A1<22> ,\DSP_PREADD_DATA.A2A1<21> ,\DSP_PREADD_DATA.A2A1<20> ,\DSP_PREADD_DATA.A2A1<19> ,\DSP_PREADD_DATA.A2A1<18> ,\DSP_PREADD_DATA.A2A1<17> ,\DSP_PREADD_DATA.A2A1<16> ,\DSP_PREADD_DATA.A2A1<15> ,\DSP_PREADD_DATA.A2A1<14> ,\DSP_PREADD_DATA.A2A1<13> ,\DSP_PREADD_DATA.A2A1<12> ,\DSP_PREADD_DATA.A2A1<11> ,\DSP_PREADD_DATA.A2A1<10> ,\DSP_PREADD_DATA.A2A1<9> ,\DSP_PREADD_DATA.A2A1<8> ,\DSP_PREADD_DATA.A2A1<7> ,\DSP_PREADD_DATA.A2A1<6> ,\DSP_PREADD_DATA.A2A1<5> ,\DSP_PREADD_DATA.A2A1<4> ,\DSP_PREADD_DATA.A2A1<3> ,\DSP_PREADD_DATA.A2A1<2> ,\DSP_PREADD_DATA.A2A1<1> ,\DSP_PREADD_DATA.A2A1<0> }),
        .AD_DATA({\DSP_PREADD_DATA.AD_DATA<26> ,\DSP_PREADD_DATA.AD_DATA<25> ,\DSP_PREADD_DATA.AD_DATA<24> ,\DSP_PREADD_DATA.AD_DATA<23> ,\DSP_PREADD_DATA.AD_DATA<22> ,\DSP_PREADD_DATA.AD_DATA<21> ,\DSP_PREADD_DATA.AD_DATA<20> ,\DSP_PREADD_DATA.AD_DATA<19> ,\DSP_PREADD_DATA.AD_DATA<18> ,\DSP_PREADD_DATA.AD_DATA<17> ,\DSP_PREADD_DATA.AD_DATA<16> ,\DSP_PREADD_DATA.AD_DATA<15> ,\DSP_PREADD_DATA.AD_DATA<14> ,\DSP_PREADD_DATA.AD_DATA<13> ,\DSP_PREADD_DATA.AD_DATA<12> ,\DSP_PREADD_DATA.AD_DATA<11> ,\DSP_PREADD_DATA.AD_DATA<10> ,\DSP_PREADD_DATA.AD_DATA<9> ,\DSP_PREADD_DATA.AD_DATA<8> ,\DSP_PREADD_DATA.AD_DATA<7> ,\DSP_PREADD_DATA.AD_DATA<6> ,\DSP_PREADD_DATA.AD_DATA<5> ,\DSP_PREADD_DATA.AD_DATA<4> ,\DSP_PREADD_DATA.AD_DATA<3> ,\DSP_PREADD_DATA.AD_DATA<2> ,\DSP_PREADD_DATA.AD_DATA<1> ,\DSP_PREADD_DATA.AD_DATA<0> }),
        .AMULT26(\DSP_MULTIPLIER.AMULT26 ),
        .B2B1({\DSP_PREADD_DATA.B2B1<17> ,\DSP_PREADD_DATA.B2B1<16> ,\DSP_PREADD_DATA.B2B1<15> ,\DSP_PREADD_DATA.B2B1<14> ,\DSP_PREADD_DATA.B2B1<13> ,\DSP_PREADD_DATA.B2B1<12> ,\DSP_PREADD_DATA.B2B1<11> ,\DSP_PREADD_DATA.B2B1<10> ,\DSP_PREADD_DATA.B2B1<9> ,\DSP_PREADD_DATA.B2B1<8> ,\DSP_PREADD_DATA.B2B1<7> ,\DSP_PREADD_DATA.B2B1<6> ,\DSP_PREADD_DATA.B2B1<5> ,\DSP_PREADD_DATA.B2B1<4> ,\DSP_PREADD_DATA.B2B1<3> ,\DSP_PREADD_DATA.B2B1<2> ,\DSP_PREADD_DATA.B2B1<1> ,\DSP_PREADD_DATA.B2B1<0> }),
        .BMULT17(\DSP_MULTIPLIER.BMULT17 ),
        .U({\DSP_MULTIPLIER.U<44> ,\DSP_MULTIPLIER.U<43> ,\DSP_MULTIPLIER.U<42> ,\DSP_MULTIPLIER.U<41> ,\DSP_MULTIPLIER.U<40> ,\DSP_MULTIPLIER.U<39> ,\DSP_MULTIPLIER.U<38> ,\DSP_MULTIPLIER.U<37> ,\DSP_MULTIPLIER.U<36> ,\DSP_MULTIPLIER.U<35> ,\DSP_MULTIPLIER.U<34> ,\DSP_MULTIPLIER.U<33> ,\DSP_MULTIPLIER.U<32> ,\DSP_MULTIPLIER.U<31> ,\DSP_MULTIPLIER.U<30> ,\DSP_MULTIPLIER.U<29> ,\DSP_MULTIPLIER.U<28> ,\DSP_MULTIPLIER.U<27> ,\DSP_MULTIPLIER.U<26> ,\DSP_MULTIPLIER.U<25> ,\DSP_MULTIPLIER.U<24> ,\DSP_MULTIPLIER.U<23> ,\DSP_MULTIPLIER.U<22> ,\DSP_MULTIPLIER.U<21> ,\DSP_MULTIPLIER.U<20> ,\DSP_MULTIPLIER.U<19> ,\DSP_MULTIPLIER.U<18> ,\DSP_MULTIPLIER.U<17> ,\DSP_MULTIPLIER.U<16> ,\DSP_MULTIPLIER.U<15> ,\DSP_MULTIPLIER.U<14> ,\DSP_MULTIPLIER.U<13> ,\DSP_MULTIPLIER.U<12> ,\DSP_MULTIPLIER.U<11> ,\DSP_MULTIPLIER.U<10> ,\DSP_MULTIPLIER.U<9> ,\DSP_MULTIPLIER.U<8> ,\DSP_MULTIPLIER.U<7> ,\DSP_MULTIPLIER.U<6> ,\DSP_MULTIPLIER.U<5> ,\DSP_MULTIPLIER.U<4> ,\DSP_MULTIPLIER.U<3> ,\DSP_MULTIPLIER.U<2> ,\DSP_MULTIPLIER.U<1> ,\DSP_MULTIPLIER.U<0> }),
        .V({\DSP_MULTIPLIER.V<44> ,\DSP_MULTIPLIER.V<43> ,\DSP_MULTIPLIER.V<42> ,\DSP_MULTIPLIER.V<41> ,\DSP_MULTIPLIER.V<40> ,\DSP_MULTIPLIER.V<39> ,\DSP_MULTIPLIER.V<38> ,\DSP_MULTIPLIER.V<37> ,\DSP_MULTIPLIER.V<36> ,\DSP_MULTIPLIER.V<35> ,\DSP_MULTIPLIER.V<34> ,\DSP_MULTIPLIER.V<33> ,\DSP_MULTIPLIER.V<32> ,\DSP_MULTIPLIER.V<31> ,\DSP_MULTIPLIER.V<30> ,\DSP_MULTIPLIER.V<29> ,\DSP_MULTIPLIER.V<28> ,\DSP_MULTIPLIER.V<27> ,\DSP_MULTIPLIER.V<26> ,\DSP_MULTIPLIER.V<25> ,\DSP_MULTIPLIER.V<24> ,\DSP_MULTIPLIER.V<23> ,\DSP_MULTIPLIER.V<22> ,\DSP_MULTIPLIER.V<21> ,\DSP_MULTIPLIER.V<20> ,\DSP_MULTIPLIER.V<19> ,\DSP_MULTIPLIER.V<18> ,\DSP_MULTIPLIER.V<17> ,\DSP_MULTIPLIER.V<16> ,\DSP_MULTIPLIER.V<15> ,\DSP_MULTIPLIER.V<14> ,\DSP_MULTIPLIER.V<13> ,\DSP_MULTIPLIER.V<12> ,\DSP_MULTIPLIER.V<11> ,\DSP_MULTIPLIER.V<10> ,\DSP_MULTIPLIER.V<9> ,\DSP_MULTIPLIER.V<8> ,\DSP_MULTIPLIER.V<7> ,\DSP_MULTIPLIER.V<6> ,\DSP_MULTIPLIER.V<5> ,\DSP_MULTIPLIER.V<4> ,\DSP_MULTIPLIER.V<3> ,\DSP_MULTIPLIER.V<2> ,\DSP_MULTIPLIER.V<1> ,\DSP_MULTIPLIER.V<0> }));
  DSP_M_DATA #(
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .MREG(0)) 
    DSP_M_DATA_INST
       (.CEM(CEM),
        .CLK(CLK),
        .RSTM(RSTM),
        .U({\DSP_MULTIPLIER.U<44> ,\DSP_MULTIPLIER.U<43> ,\DSP_MULTIPLIER.U<42> ,\DSP_MULTIPLIER.U<41> ,\DSP_MULTIPLIER.U<40> ,\DSP_MULTIPLIER.U<39> ,\DSP_MULTIPLIER.U<38> ,\DSP_MULTIPLIER.U<37> ,\DSP_MULTIPLIER.U<36> ,\DSP_MULTIPLIER.U<35> ,\DSP_MULTIPLIER.U<34> ,\DSP_MULTIPLIER.U<33> ,\DSP_MULTIPLIER.U<32> ,\DSP_MULTIPLIER.U<31> ,\DSP_MULTIPLIER.U<30> ,\DSP_MULTIPLIER.U<29> ,\DSP_MULTIPLIER.U<28> ,\DSP_MULTIPLIER.U<27> ,\DSP_MULTIPLIER.U<26> ,\DSP_MULTIPLIER.U<25> ,\DSP_MULTIPLIER.U<24> ,\DSP_MULTIPLIER.U<23> ,\DSP_MULTIPLIER.U<22> ,\DSP_MULTIPLIER.U<21> ,\DSP_MULTIPLIER.U<20> ,\DSP_MULTIPLIER.U<19> ,\DSP_MULTIPLIER.U<18> ,\DSP_MULTIPLIER.U<17> ,\DSP_MULTIPLIER.U<16> ,\DSP_MULTIPLIER.U<15> ,\DSP_MULTIPLIER.U<14> ,\DSP_MULTIPLIER.U<13> ,\DSP_MULTIPLIER.U<12> ,\DSP_MULTIPLIER.U<11> ,\DSP_MULTIPLIER.U<10> ,\DSP_MULTIPLIER.U<9> ,\DSP_MULTIPLIER.U<8> ,\DSP_MULTIPLIER.U<7> ,\DSP_MULTIPLIER.U<6> ,\DSP_MULTIPLIER.U<5> ,\DSP_MULTIPLIER.U<4> ,\DSP_MULTIPLIER.U<3> ,\DSP_MULTIPLIER.U<2> ,\DSP_MULTIPLIER.U<1> ,\DSP_MULTIPLIER.U<0> }),
        .U_DATA({\DSP_M_DATA.U_DATA<44> ,\DSP_M_DATA.U_DATA<43> ,\DSP_M_DATA.U_DATA<42> ,\DSP_M_DATA.U_DATA<41> ,\DSP_M_DATA.U_DATA<40> ,\DSP_M_DATA.U_DATA<39> ,\DSP_M_DATA.U_DATA<38> ,\DSP_M_DATA.U_DATA<37> ,\DSP_M_DATA.U_DATA<36> ,\DSP_M_DATA.U_DATA<35> ,\DSP_M_DATA.U_DATA<34> ,\DSP_M_DATA.U_DATA<33> ,\DSP_M_DATA.U_DATA<32> ,\DSP_M_DATA.U_DATA<31> ,\DSP_M_DATA.U_DATA<30> ,\DSP_M_DATA.U_DATA<29> ,\DSP_M_DATA.U_DATA<28> ,\DSP_M_DATA.U_DATA<27> ,\DSP_M_DATA.U_DATA<26> ,\DSP_M_DATA.U_DATA<25> ,\DSP_M_DATA.U_DATA<24> ,\DSP_M_DATA.U_DATA<23> ,\DSP_M_DATA.U_DATA<22> ,\DSP_M_DATA.U_DATA<21> ,\DSP_M_DATA.U_DATA<20> ,\DSP_M_DATA.U_DATA<19> ,\DSP_M_DATA.U_DATA<18> ,\DSP_M_DATA.U_DATA<17> ,\DSP_M_DATA.U_DATA<16> ,\DSP_M_DATA.U_DATA<15> ,\DSP_M_DATA.U_DATA<14> ,\DSP_M_DATA.U_DATA<13> ,\DSP_M_DATA.U_DATA<12> ,\DSP_M_DATA.U_DATA<11> ,\DSP_M_DATA.U_DATA<10> ,\DSP_M_DATA.U_DATA<9> ,\DSP_M_DATA.U_DATA<8> ,\DSP_M_DATA.U_DATA<7> ,\DSP_M_DATA.U_DATA<6> ,\DSP_M_DATA.U_DATA<5> ,\DSP_M_DATA.U_DATA<4> ,\DSP_M_DATA.U_DATA<3> ,\DSP_M_DATA.U_DATA<2> ,\DSP_M_DATA.U_DATA<1> ,\DSP_M_DATA.U_DATA<0> }),
        .V({\DSP_MULTIPLIER.V<44> ,\DSP_MULTIPLIER.V<43> ,\DSP_MULTIPLIER.V<42> ,\DSP_MULTIPLIER.V<41> ,\DSP_MULTIPLIER.V<40> ,\DSP_MULTIPLIER.V<39> ,\DSP_MULTIPLIER.V<38> ,\DSP_MULTIPLIER.V<37> ,\DSP_MULTIPLIER.V<36> ,\DSP_MULTIPLIER.V<35> ,\DSP_MULTIPLIER.V<34> ,\DSP_MULTIPLIER.V<33> ,\DSP_MULTIPLIER.V<32> ,\DSP_MULTIPLIER.V<31> ,\DSP_MULTIPLIER.V<30> ,\DSP_MULTIPLIER.V<29> ,\DSP_MULTIPLIER.V<28> ,\DSP_MULTIPLIER.V<27> ,\DSP_MULTIPLIER.V<26> ,\DSP_MULTIPLIER.V<25> ,\DSP_MULTIPLIER.V<24> ,\DSP_MULTIPLIER.V<23> ,\DSP_MULTIPLIER.V<22> ,\DSP_MULTIPLIER.V<21> ,\DSP_MULTIPLIER.V<20> ,\DSP_MULTIPLIER.V<19> ,\DSP_MULTIPLIER.V<18> ,\DSP_MULTIPLIER.V<17> ,\DSP_MULTIPLIER.V<16> ,\DSP_MULTIPLIER.V<15> ,\DSP_MULTIPLIER.V<14> ,\DSP_MULTIPLIER.V<13> ,\DSP_MULTIPLIER.V<12> ,\DSP_MULTIPLIER.V<11> ,\DSP_MULTIPLIER.V<10> ,\DSP_MULTIPLIER.V<9> ,\DSP_MULTIPLIER.V<8> ,\DSP_MULTIPLIER.V<7> ,\DSP_MULTIPLIER.V<6> ,\DSP_MULTIPLIER.V<5> ,\DSP_MULTIPLIER.V<4> ,\DSP_MULTIPLIER.V<3> ,\DSP_MULTIPLIER.V<2> ,\DSP_MULTIPLIER.V<1> ,\DSP_MULTIPLIER.V<0> }),
        .V_DATA({\DSP_M_DATA.V_DATA<44> ,\DSP_M_DATA.V_DATA<43> ,\DSP_M_DATA.V_DATA<42> ,\DSP_M_DATA.V_DATA<41> ,\DSP_M_DATA.V_DATA<40> ,\DSP_M_DATA.V_DATA<39> ,\DSP_M_DATA.V_DATA<38> ,\DSP_M_DATA.V_DATA<37> ,\DSP_M_DATA.V_DATA<36> ,\DSP_M_DATA.V_DATA<35> ,\DSP_M_DATA.V_DATA<34> ,\DSP_M_DATA.V_DATA<33> ,\DSP_M_DATA.V_DATA<32> ,\DSP_M_DATA.V_DATA<31> ,\DSP_M_DATA.V_DATA<30> ,\DSP_M_DATA.V_DATA<29> ,\DSP_M_DATA.V_DATA<28> ,\DSP_M_DATA.V_DATA<27> ,\DSP_M_DATA.V_DATA<26> ,\DSP_M_DATA.V_DATA<25> ,\DSP_M_DATA.V_DATA<24> ,\DSP_M_DATA.V_DATA<23> ,\DSP_M_DATA.V_DATA<22> ,\DSP_M_DATA.V_DATA<21> ,\DSP_M_DATA.V_DATA<20> ,\DSP_M_DATA.V_DATA<19> ,\DSP_M_DATA.V_DATA<18> ,\DSP_M_DATA.V_DATA<17> ,\DSP_M_DATA.V_DATA<16> ,\DSP_M_DATA.V_DATA<15> ,\DSP_M_DATA.V_DATA<14> ,\DSP_M_DATA.V_DATA<13> ,\DSP_M_DATA.V_DATA<12> ,\DSP_M_DATA.V_DATA<11> ,\DSP_M_DATA.V_DATA<10> ,\DSP_M_DATA.V_DATA<9> ,\DSP_M_DATA.V_DATA<8> ,\DSP_M_DATA.V_DATA<7> ,\DSP_M_DATA.V_DATA<6> ,\DSP_M_DATA.V_DATA<5> ,\DSP_M_DATA.V_DATA<4> ,\DSP_M_DATA.V_DATA<3> ,\DSP_M_DATA.V_DATA<2> ,\DSP_M_DATA.V_DATA<1> ,\DSP_M_DATA.V_DATA<0> }));
  DSP_OUTPUT #(
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h3FFFFFFFFFFF),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_PATTERN_DETECT("NO_PATDET")) 
    DSP_OUTPUT_INST
       (.ALUMODE10(\DSP_ALU.ALUMODE10 ),
        .ALU_OUT({\DSP_ALU.ALU_OUT<47> ,\DSP_ALU.ALU_OUT<46> ,\DSP_ALU.ALU_OUT<45> ,\DSP_ALU.ALU_OUT<44> ,\DSP_ALU.ALU_OUT<43> ,\DSP_ALU.ALU_OUT<42> ,\DSP_ALU.ALU_OUT<41> ,\DSP_ALU.ALU_OUT<40> ,\DSP_ALU.ALU_OUT<39> ,\DSP_ALU.ALU_OUT<38> ,\DSP_ALU.ALU_OUT<37> ,\DSP_ALU.ALU_OUT<36> ,\DSP_ALU.ALU_OUT<35> ,\DSP_ALU.ALU_OUT<34> ,\DSP_ALU.ALU_OUT<33> ,\DSP_ALU.ALU_OUT<32> ,\DSP_ALU.ALU_OUT<31> ,\DSP_ALU.ALU_OUT<30> ,\DSP_ALU.ALU_OUT<29> ,\DSP_ALU.ALU_OUT<28> ,\DSP_ALU.ALU_OUT<27> ,\DSP_ALU.ALU_OUT<26> ,\DSP_ALU.ALU_OUT<25> ,\DSP_ALU.ALU_OUT<24> ,\DSP_ALU.ALU_OUT<23> ,\DSP_ALU.ALU_OUT<22> ,\DSP_ALU.ALU_OUT<21> ,\DSP_ALU.ALU_OUT<20> ,\DSP_ALU.ALU_OUT<19> ,\DSP_ALU.ALU_OUT<18> ,\DSP_ALU.ALU_OUT<17> ,\DSP_ALU.ALU_OUT<16> ,\DSP_ALU.ALU_OUT<15> ,\DSP_ALU.ALU_OUT<14> ,\DSP_ALU.ALU_OUT<13> ,\DSP_ALU.ALU_OUT<12> ,\DSP_ALU.ALU_OUT<11> ,\DSP_ALU.ALU_OUT<10> ,\DSP_ALU.ALU_OUT<9> ,\DSP_ALU.ALU_OUT<8> ,\DSP_ALU.ALU_OUT<7> ,\DSP_ALU.ALU_OUT<6> ,\DSP_ALU.ALU_OUT<5> ,\DSP_ALU.ALU_OUT<4> ,\DSP_ALU.ALU_OUT<3> ,\DSP_ALU.ALU_OUT<2> ,\DSP_ALU.ALU_OUT<1> ,\DSP_ALU.ALU_OUT<0> }),
        .CARRYCASCOUT(CARRYCASCOUT),
        .CARRYOUT({\CARRYOUT[3] ,\CARRYOUT[2] ,\CARRYOUT[1] ,\CARRYOUT[0] }),
        .CCOUT_FB(\DSP_OUTPUT.CCOUT_FB ),
        .CEP(CEP),
        .CLK(CLK),
        .COUT({\DSP_ALU.COUT<3> ,\DSP_ALU.COUT<2> ,\DSP_ALU.COUT<1> ,\DSP_ALU.COUT<0> }),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .MULTSIGNOUT(MULTSIGNOUT),
        .MULTSIGN_ALU(\DSP_ALU.MULTSIGN_ALU ),
        .OVERFLOW(OVERFLOW),
        .P({\P[47] ,\P[46] ,\P[45] ,\P[44] ,\P[43] ,\P[42] ,\P[41] ,\P[40] ,\P[39] ,\P[38] ,\P[37] ,\P[36] ,\P[35] ,\P[34] ,\P[33] ,\P[32] ,\P[31] ,\P[30] ,\P[29] ,\P[28] ,\P[27] ,\P[26] ,\P[25] ,\P[24] ,\P[23] ,\P[22] ,\P[21] ,\P[20] ,\P[19] ,\P[18] ,\P[17] ,\P[16] ,\P[15] ,\P[14] ,\P[13] ,\P[12] ,\P[11] ,\P[10] ,\P[9] ,\P[8] ,\P[7] ,\P[6] ,\P[5] ,\P[4] ,\P[3] ,\P[2] ,\P[1] ,\P[0] }),
        .PATTERN_B_DETECT(PATTERNBDETECT),
        .PATTERN_DETECT(PATTERNDETECT),
        .PCOUT({\PCOUT[47] ,\PCOUT[46] ,\PCOUT[45] ,\PCOUT[44] ,\PCOUT[43] ,\PCOUT[42] ,\PCOUT[41] ,\PCOUT[40] ,\PCOUT[39] ,\PCOUT[38] ,\PCOUT[37] ,\PCOUT[36] ,\PCOUT[35] ,\PCOUT[34] ,\PCOUT[33] ,\PCOUT[32] ,\PCOUT[31] ,\PCOUT[30] ,\PCOUT[29] ,\PCOUT[28] ,\PCOUT[27] ,\PCOUT[26] ,\PCOUT[25] ,\PCOUT[24] ,\PCOUT[23] ,\PCOUT[22] ,\PCOUT[21] ,\PCOUT[20] ,\PCOUT[19] ,\PCOUT[18] ,\PCOUT[17] ,\PCOUT[16] ,\PCOUT[15] ,\PCOUT[14] ,\PCOUT[13] ,\PCOUT[12] ,\PCOUT[11] ,\PCOUT[10] ,\PCOUT[9] ,\PCOUT[8] ,\PCOUT[7] ,\PCOUT[6] ,\PCOUT[5] ,\PCOUT[4] ,\PCOUT[3] ,\PCOUT[2] ,\PCOUT[1] ,\PCOUT[0] }),
        .P_FDBK({\DSP_OUTPUT.P_FDBK<47> ,\DSP_OUTPUT.P_FDBK<46> ,\DSP_OUTPUT.P_FDBK<45> ,\DSP_OUTPUT.P_FDBK<44> ,\DSP_OUTPUT.P_FDBK<43> ,\DSP_OUTPUT.P_FDBK<42> ,\DSP_OUTPUT.P_FDBK<41> ,\DSP_OUTPUT.P_FDBK<40> ,\DSP_OUTPUT.P_FDBK<39> ,\DSP_OUTPUT.P_FDBK<38> ,\DSP_OUTPUT.P_FDBK<37> ,\DSP_OUTPUT.P_FDBK<36> ,\DSP_OUTPUT.P_FDBK<35> ,\DSP_OUTPUT.P_FDBK<34> ,\DSP_OUTPUT.P_FDBK<33> ,\DSP_OUTPUT.P_FDBK<32> ,\DSP_OUTPUT.P_FDBK<31> ,\DSP_OUTPUT.P_FDBK<30> ,\DSP_OUTPUT.P_FDBK<29> ,\DSP_OUTPUT.P_FDBK<28> ,\DSP_OUTPUT.P_FDBK<27> ,\DSP_OUTPUT.P_FDBK<26> ,\DSP_OUTPUT.P_FDBK<25> ,\DSP_OUTPUT.P_FDBK<24> ,\DSP_OUTPUT.P_FDBK<23> ,\DSP_OUTPUT.P_FDBK<22> ,\DSP_OUTPUT.P_FDBK<21> ,\DSP_OUTPUT.P_FDBK<20> ,\DSP_OUTPUT.P_FDBK<19> ,\DSP_OUTPUT.P_FDBK<18> ,\DSP_OUTPUT.P_FDBK<17> ,\DSP_OUTPUT.P_FDBK<16> ,\DSP_OUTPUT.P_FDBK<15> ,\DSP_OUTPUT.P_FDBK<14> ,\DSP_OUTPUT.P_FDBK<13> ,\DSP_OUTPUT.P_FDBK<12> ,\DSP_OUTPUT.P_FDBK<11> ,\DSP_OUTPUT.P_FDBK<10> ,\DSP_OUTPUT.P_FDBK<9> ,\DSP_OUTPUT.P_FDBK<8> ,\DSP_OUTPUT.P_FDBK<7> ,\DSP_OUTPUT.P_FDBK<6> ,\DSP_OUTPUT.P_FDBK<5> ,\DSP_OUTPUT.P_FDBK<4> ,\DSP_OUTPUT.P_FDBK<3> ,\DSP_OUTPUT.P_FDBK<2> ,\DSP_OUTPUT.P_FDBK<1> ,\DSP_OUTPUT.P_FDBK<0> }),
        .P_FDBK_47(\DSP_OUTPUT.P_FDBK_47 ),
        .RSTP(RSTP),
        .UNDERFLOW(UNDERFLOW),
        .XOROUT({\XOROUT[7] ,\XOROUT[6] ,\XOROUT[5] ,\XOROUT[4] ,\XOROUT[3] ,\XOROUT[2] ,\XOROUT[1] ,\XOROUT[0] }),
        .XOR_MX({\DSP_ALU.XOR_MX<7> ,\DSP_ALU.XOR_MX<6> ,\DSP_ALU.XOR_MX<5> ,\DSP_ALU.XOR_MX<4> ,\DSP_ALU.XOR_MX<3> ,\DSP_ALU.XOR_MX<2> ,\DSP_ALU.XOR_MX<1> ,\DSP_ALU.XOR_MX<0> }));
  DSP_PREADD_DATA #(
    .ADREG(1),
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .DREG(1),
    .INMODEREG(0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .PREADDINSEL("A"),
    .USE_MULT("MULTIPLY")) 
    DSP_PREADD_DATA_INST
       (.A1_DATA({\DSP_A_B_DATA.A1_DATA<26> ,\DSP_A_B_DATA.A1_DATA<25> ,\DSP_A_B_DATA.A1_DATA<24> ,\DSP_A_B_DATA.A1_DATA<23> ,\DSP_A_B_DATA.A1_DATA<22> ,\DSP_A_B_DATA.A1_DATA<21> ,\DSP_A_B_DATA.A1_DATA<20> ,\DSP_A_B_DATA.A1_DATA<19> ,\DSP_A_B_DATA.A1_DATA<18> ,\DSP_A_B_DATA.A1_DATA<17> ,\DSP_A_B_DATA.A1_DATA<16> ,\DSP_A_B_DATA.A1_DATA<15> ,\DSP_A_B_DATA.A1_DATA<14> ,\DSP_A_B_DATA.A1_DATA<13> ,\DSP_A_B_DATA.A1_DATA<12> ,\DSP_A_B_DATA.A1_DATA<11> ,\DSP_A_B_DATA.A1_DATA<10> ,\DSP_A_B_DATA.A1_DATA<9> ,\DSP_A_B_DATA.A1_DATA<8> ,\DSP_A_B_DATA.A1_DATA<7> ,\DSP_A_B_DATA.A1_DATA<6> ,\DSP_A_B_DATA.A1_DATA<5> ,\DSP_A_B_DATA.A1_DATA<4> ,\DSP_A_B_DATA.A1_DATA<3> ,\DSP_A_B_DATA.A1_DATA<2> ,\DSP_A_B_DATA.A1_DATA<1> ,\DSP_A_B_DATA.A1_DATA<0> }),
        .A2A1({\DSP_PREADD_DATA.A2A1<26> ,\DSP_PREADD_DATA.A2A1<25> ,\DSP_PREADD_DATA.A2A1<24> ,\DSP_PREADD_DATA.A2A1<23> ,\DSP_PREADD_DATA.A2A1<22> ,\DSP_PREADD_DATA.A2A1<21> ,\DSP_PREADD_DATA.A2A1<20> ,\DSP_PREADD_DATA.A2A1<19> ,\DSP_PREADD_DATA.A2A1<18> ,\DSP_PREADD_DATA.A2A1<17> ,\DSP_PREADD_DATA.A2A1<16> ,\DSP_PREADD_DATA.A2A1<15> ,\DSP_PREADD_DATA.A2A1<14> ,\DSP_PREADD_DATA.A2A1<13> ,\DSP_PREADD_DATA.A2A1<12> ,\DSP_PREADD_DATA.A2A1<11> ,\DSP_PREADD_DATA.A2A1<10> ,\DSP_PREADD_DATA.A2A1<9> ,\DSP_PREADD_DATA.A2A1<8> ,\DSP_PREADD_DATA.A2A1<7> ,\DSP_PREADD_DATA.A2A1<6> ,\DSP_PREADD_DATA.A2A1<5> ,\DSP_PREADD_DATA.A2A1<4> ,\DSP_PREADD_DATA.A2A1<3> ,\DSP_PREADD_DATA.A2A1<2> ,\DSP_PREADD_DATA.A2A1<1> ,\DSP_PREADD_DATA.A2A1<0> }),
        .A2_DATA({\DSP_A_B_DATA.A2_DATA<26> ,\DSP_A_B_DATA.A2_DATA<25> ,\DSP_A_B_DATA.A2_DATA<24> ,\DSP_A_B_DATA.A2_DATA<23> ,\DSP_A_B_DATA.A2_DATA<22> ,\DSP_A_B_DATA.A2_DATA<21> ,\DSP_A_B_DATA.A2_DATA<20> ,\DSP_A_B_DATA.A2_DATA<19> ,\DSP_A_B_DATA.A2_DATA<18> ,\DSP_A_B_DATA.A2_DATA<17> ,\DSP_A_B_DATA.A2_DATA<16> ,\DSP_A_B_DATA.A2_DATA<15> ,\DSP_A_B_DATA.A2_DATA<14> ,\DSP_A_B_DATA.A2_DATA<13> ,\DSP_A_B_DATA.A2_DATA<12> ,\DSP_A_B_DATA.A2_DATA<11> ,\DSP_A_B_DATA.A2_DATA<10> ,\DSP_A_B_DATA.A2_DATA<9> ,\DSP_A_B_DATA.A2_DATA<8> ,\DSP_A_B_DATA.A2_DATA<7> ,\DSP_A_B_DATA.A2_DATA<6> ,\DSP_A_B_DATA.A2_DATA<5> ,\DSP_A_B_DATA.A2_DATA<4> ,\DSP_A_B_DATA.A2_DATA<3> ,\DSP_A_B_DATA.A2_DATA<2> ,\DSP_A_B_DATA.A2_DATA<1> ,\DSP_A_B_DATA.A2_DATA<0> }),
        .AD({\DSP_PREADD.AD<26> ,\DSP_PREADD.AD<25> ,\DSP_PREADD.AD<24> ,\DSP_PREADD.AD<23> ,\DSP_PREADD.AD<22> ,\DSP_PREADD.AD<21> ,\DSP_PREADD.AD<20> ,\DSP_PREADD.AD<19> ,\DSP_PREADD.AD<18> ,\DSP_PREADD.AD<17> ,\DSP_PREADD.AD<16> ,\DSP_PREADD.AD<15> ,\DSP_PREADD.AD<14> ,\DSP_PREADD.AD<13> ,\DSP_PREADD.AD<12> ,\DSP_PREADD.AD<11> ,\DSP_PREADD.AD<10> ,\DSP_PREADD.AD<9> ,\DSP_PREADD.AD<8> ,\DSP_PREADD.AD<7> ,\DSP_PREADD.AD<6> ,\DSP_PREADD.AD<5> ,\DSP_PREADD.AD<4> ,\DSP_PREADD.AD<3> ,\DSP_PREADD.AD<2> ,\DSP_PREADD.AD<1> ,\DSP_PREADD.AD<0> }),
        .ADDSUB(\DSP_PREADD_DATA.ADDSUB ),
        .AD_DATA({\DSP_PREADD_DATA.AD_DATA<26> ,\DSP_PREADD_DATA.AD_DATA<25> ,\DSP_PREADD_DATA.AD_DATA<24> ,\DSP_PREADD_DATA.AD_DATA<23> ,\DSP_PREADD_DATA.AD_DATA<22> ,\DSP_PREADD_DATA.AD_DATA<21> ,\DSP_PREADD_DATA.AD_DATA<20> ,\DSP_PREADD_DATA.AD_DATA<19> ,\DSP_PREADD_DATA.AD_DATA<18> ,\DSP_PREADD_DATA.AD_DATA<17> ,\DSP_PREADD_DATA.AD_DATA<16> ,\DSP_PREADD_DATA.AD_DATA<15> ,\DSP_PREADD_DATA.AD_DATA<14> ,\DSP_PREADD_DATA.AD_DATA<13> ,\DSP_PREADD_DATA.AD_DATA<12> ,\DSP_PREADD_DATA.AD_DATA<11> ,\DSP_PREADD_DATA.AD_DATA<10> ,\DSP_PREADD_DATA.AD_DATA<9> ,\DSP_PREADD_DATA.AD_DATA<8> ,\DSP_PREADD_DATA.AD_DATA<7> ,\DSP_PREADD_DATA.AD_DATA<6> ,\DSP_PREADD_DATA.AD_DATA<5> ,\DSP_PREADD_DATA.AD_DATA<4> ,\DSP_PREADD_DATA.AD_DATA<3> ,\DSP_PREADD_DATA.AD_DATA<2> ,\DSP_PREADD_DATA.AD_DATA<1> ,\DSP_PREADD_DATA.AD_DATA<0> }),
        .B1_DATA({\DSP_A_B_DATA.B1_DATA<17> ,\DSP_A_B_DATA.B1_DATA<16> ,\DSP_A_B_DATA.B1_DATA<15> ,\DSP_A_B_DATA.B1_DATA<14> ,\DSP_A_B_DATA.B1_DATA<13> ,\DSP_A_B_DATA.B1_DATA<12> ,\DSP_A_B_DATA.B1_DATA<11> ,\DSP_A_B_DATA.B1_DATA<10> ,\DSP_A_B_DATA.B1_DATA<9> ,\DSP_A_B_DATA.B1_DATA<8> ,\DSP_A_B_DATA.B1_DATA<7> ,\DSP_A_B_DATA.B1_DATA<6> ,\DSP_A_B_DATA.B1_DATA<5> ,\DSP_A_B_DATA.B1_DATA<4> ,\DSP_A_B_DATA.B1_DATA<3> ,\DSP_A_B_DATA.B1_DATA<2> ,\DSP_A_B_DATA.B1_DATA<1> ,\DSP_A_B_DATA.B1_DATA<0> }),
        .B2B1({\DSP_PREADD_DATA.B2B1<17> ,\DSP_PREADD_DATA.B2B1<16> ,\DSP_PREADD_DATA.B2B1<15> ,\DSP_PREADD_DATA.B2B1<14> ,\DSP_PREADD_DATA.B2B1<13> ,\DSP_PREADD_DATA.B2B1<12> ,\DSP_PREADD_DATA.B2B1<11> ,\DSP_PREADD_DATA.B2B1<10> ,\DSP_PREADD_DATA.B2B1<9> ,\DSP_PREADD_DATA.B2B1<8> ,\DSP_PREADD_DATA.B2B1<7> ,\DSP_PREADD_DATA.B2B1<6> ,\DSP_PREADD_DATA.B2B1<5> ,\DSP_PREADD_DATA.B2B1<4> ,\DSP_PREADD_DATA.B2B1<3> ,\DSP_PREADD_DATA.B2B1<2> ,\DSP_PREADD_DATA.B2B1<1> ,\DSP_PREADD_DATA.B2B1<0> }),
        .B2_DATA({\DSP_A_B_DATA.B2_DATA<17> ,\DSP_A_B_DATA.B2_DATA<16> ,\DSP_A_B_DATA.B2_DATA<15> ,\DSP_A_B_DATA.B2_DATA<14> ,\DSP_A_B_DATA.B2_DATA<13> ,\DSP_A_B_DATA.B2_DATA<12> ,\DSP_A_B_DATA.B2_DATA<11> ,\DSP_A_B_DATA.B2_DATA<10> ,\DSP_A_B_DATA.B2_DATA<9> ,\DSP_A_B_DATA.B2_DATA<8> ,\DSP_A_B_DATA.B2_DATA<7> ,\DSP_A_B_DATA.B2_DATA<6> ,\DSP_A_B_DATA.B2_DATA<5> ,\DSP_A_B_DATA.B2_DATA<4> ,\DSP_A_B_DATA.B2_DATA<3> ,\DSP_A_B_DATA.B2_DATA<2> ,\DSP_A_B_DATA.B2_DATA<1> ,\DSP_A_B_DATA.B2_DATA<0> }),
        .CEAD(CEAD),
        .CED(CED),
        .CEINMODE(CEINMODE),
        .CLK(CLK),
        .DIN({\D[26] ,\D[25] ,\D[24] ,\D[23] ,\D[22] ,\D[21] ,\D[20] ,\D[19] ,\D[18] ,\D[17] ,\D[16] ,\D[15] ,\D[14] ,\D[13] ,\D[12] ,\D[11] ,\D[10] ,\D[9] ,\D[8] ,\D[7] ,\D[6] ,\D[5] ,\D[4] ,\D[3] ,\D[2] ,\D[1] ,\D[0] }),
        .D_DATA({\DSP_PREADD_DATA.D_DATA<26> ,\DSP_PREADD_DATA.D_DATA<25> ,\DSP_PREADD_DATA.D_DATA<24> ,\DSP_PREADD_DATA.D_DATA<23> ,\DSP_PREADD_DATA.D_DATA<22> ,\DSP_PREADD_DATA.D_DATA<21> ,\DSP_PREADD_DATA.D_DATA<20> ,\DSP_PREADD_DATA.D_DATA<19> ,\DSP_PREADD_DATA.D_DATA<18> ,\DSP_PREADD_DATA.D_DATA<17> ,\DSP_PREADD_DATA.D_DATA<16> ,\DSP_PREADD_DATA.D_DATA<15> ,\DSP_PREADD_DATA.D_DATA<14> ,\DSP_PREADD_DATA.D_DATA<13> ,\DSP_PREADD_DATA.D_DATA<12> ,\DSP_PREADD_DATA.D_DATA<11> ,\DSP_PREADD_DATA.D_DATA<10> ,\DSP_PREADD_DATA.D_DATA<9> ,\DSP_PREADD_DATA.D_DATA<8> ,\DSP_PREADD_DATA.D_DATA<7> ,\DSP_PREADD_DATA.D_DATA<6> ,\DSP_PREADD_DATA.D_DATA<5> ,\DSP_PREADD_DATA.D_DATA<4> ,\DSP_PREADD_DATA.D_DATA<3> ,\DSP_PREADD_DATA.D_DATA<2> ,\DSP_PREADD_DATA.D_DATA<1> ,\DSP_PREADD_DATA.D_DATA<0> }),
        .INMODE({\INMODE[4] ,\INMODE[3] ,\INMODE[2] ,\INMODE[1] ,\INMODE[0] }),
        .INMODE_2(\DSP_PREADD_DATA.INMODE_2 ),
        .PREADD_AB({\DSP_PREADD_DATA.PREADD_AB<26> ,\DSP_PREADD_DATA.PREADD_AB<25> ,\DSP_PREADD_DATA.PREADD_AB<24> ,\DSP_PREADD_DATA.PREADD_AB<23> ,\DSP_PREADD_DATA.PREADD_AB<22> ,\DSP_PREADD_DATA.PREADD_AB<21> ,\DSP_PREADD_DATA.PREADD_AB<20> ,\DSP_PREADD_DATA.PREADD_AB<19> ,\DSP_PREADD_DATA.PREADD_AB<18> ,\DSP_PREADD_DATA.PREADD_AB<17> ,\DSP_PREADD_DATA.PREADD_AB<16> ,\DSP_PREADD_DATA.PREADD_AB<15> ,\DSP_PREADD_DATA.PREADD_AB<14> ,\DSP_PREADD_DATA.PREADD_AB<13> ,\DSP_PREADD_DATA.PREADD_AB<12> ,\DSP_PREADD_DATA.PREADD_AB<11> ,\DSP_PREADD_DATA.PREADD_AB<10> ,\DSP_PREADD_DATA.PREADD_AB<9> ,\DSP_PREADD_DATA.PREADD_AB<8> ,\DSP_PREADD_DATA.PREADD_AB<7> ,\DSP_PREADD_DATA.PREADD_AB<6> ,\DSP_PREADD_DATA.PREADD_AB<5> ,\DSP_PREADD_DATA.PREADD_AB<4> ,\DSP_PREADD_DATA.PREADD_AB<3> ,\DSP_PREADD_DATA.PREADD_AB<2> ,\DSP_PREADD_DATA.PREADD_AB<1> ,\DSP_PREADD_DATA.PREADD_AB<0> }),
        .RSTD(RSTD),
        .RSTINMODE(RSTINMODE));
  DSP_PREADD DSP_PREADD_INST
       (.AD({\DSP_PREADD.AD<26> ,\DSP_PREADD.AD<25> ,\DSP_PREADD.AD<24> ,\DSP_PREADD.AD<23> ,\DSP_PREADD.AD<22> ,\DSP_PREADD.AD<21> ,\DSP_PREADD.AD<20> ,\DSP_PREADD.AD<19> ,\DSP_PREADD.AD<18> ,\DSP_PREADD.AD<17> ,\DSP_PREADD.AD<16> ,\DSP_PREADD.AD<15> ,\DSP_PREADD.AD<14> ,\DSP_PREADD.AD<13> ,\DSP_PREADD.AD<12> ,\DSP_PREADD.AD<11> ,\DSP_PREADD.AD<10> ,\DSP_PREADD.AD<9> ,\DSP_PREADD.AD<8> ,\DSP_PREADD.AD<7> ,\DSP_PREADD.AD<6> ,\DSP_PREADD.AD<5> ,\DSP_PREADD.AD<4> ,\DSP_PREADD.AD<3> ,\DSP_PREADD.AD<2> ,\DSP_PREADD.AD<1> ,\DSP_PREADD.AD<0> }),
        .ADDSUB(\DSP_PREADD_DATA.ADDSUB ),
        .D_DATA({\DSP_PREADD_DATA.D_DATA<26> ,\DSP_PREADD_DATA.D_DATA<25> ,\DSP_PREADD_DATA.D_DATA<24> ,\DSP_PREADD_DATA.D_DATA<23> ,\DSP_PREADD_DATA.D_DATA<22> ,\DSP_PREADD_DATA.D_DATA<21> ,\DSP_PREADD_DATA.D_DATA<20> ,\DSP_PREADD_DATA.D_DATA<19> ,\DSP_PREADD_DATA.D_DATA<18> ,\DSP_PREADD_DATA.D_DATA<17> ,\DSP_PREADD_DATA.D_DATA<16> ,\DSP_PREADD_DATA.D_DATA<15> ,\DSP_PREADD_DATA.D_DATA<14> ,\DSP_PREADD_DATA.D_DATA<13> ,\DSP_PREADD_DATA.D_DATA<12> ,\DSP_PREADD_DATA.D_DATA<11> ,\DSP_PREADD_DATA.D_DATA<10> ,\DSP_PREADD_DATA.D_DATA<9> ,\DSP_PREADD_DATA.D_DATA<8> ,\DSP_PREADD_DATA.D_DATA<7> ,\DSP_PREADD_DATA.D_DATA<6> ,\DSP_PREADD_DATA.D_DATA<5> ,\DSP_PREADD_DATA.D_DATA<4> ,\DSP_PREADD_DATA.D_DATA<3> ,\DSP_PREADD_DATA.D_DATA<2> ,\DSP_PREADD_DATA.D_DATA<1> ,\DSP_PREADD_DATA.D_DATA<0> }),
        .INMODE2(\DSP_PREADD_DATA.INMODE_2 ),
        .PREADD_AB({\DSP_PREADD_DATA.PREADD_AB<26> ,\DSP_PREADD_DATA.PREADD_AB<25> ,\DSP_PREADD_DATA.PREADD_AB<24> ,\DSP_PREADD_DATA.PREADD_AB<23> ,\DSP_PREADD_DATA.PREADD_AB<22> ,\DSP_PREADD_DATA.PREADD_AB<21> ,\DSP_PREADD_DATA.PREADD_AB<20> ,\DSP_PREADD_DATA.PREADD_AB<19> ,\DSP_PREADD_DATA.PREADD_AB<18> ,\DSP_PREADD_DATA.PREADD_AB<17> ,\DSP_PREADD_DATA.PREADD_AB<16> ,\DSP_PREADD_DATA.PREADD_AB<15> ,\DSP_PREADD_DATA.PREADD_AB<14> ,\DSP_PREADD_DATA.PREADD_AB<13> ,\DSP_PREADD_DATA.PREADD_AB<12> ,\DSP_PREADD_DATA.PREADD_AB<11> ,\DSP_PREADD_DATA.PREADD_AB<10> ,\DSP_PREADD_DATA.PREADD_AB<9> ,\DSP_PREADD_DATA.PREADD_AB<8> ,\DSP_PREADD_DATA.PREADD_AB<7> ,\DSP_PREADD_DATA.PREADD_AB<6> ,\DSP_PREADD_DATA.PREADD_AB<5> ,\DSP_PREADD_DATA.PREADD_AB<4> ,\DSP_PREADD_DATA.PREADD_AB<3> ,\DSP_PREADD_DATA.PREADD_AB<2> ,\DSP_PREADD_DATA.PREADD_AB<1> ,\DSP_PREADD_DATA.PREADD_AB<0> }));
endmodule

module DSP48E2_HD32740
   (ACOUT,
    BCOUT,
    CARRYCASCOUT,
    CARRYOUT,
    MULTSIGNOUT,
    OVERFLOW,
    PATTERNBDETECT,
    PATTERNDETECT,
    PCOUT,
    P,
    UNDERFLOW,
    XOROUT,
    ACIN,
    ALUMODE,
    A,
    BCIN,
    B,
    CARRYCASCIN,
    CARRYIN,
    CARRYINSEL,
    CEA1,
    CEA2,
    CEAD,
    CEALUMODE,
    CEB1,
    CEB2,
    CEC,
    CECARRYIN,
    CECTRL,
    CED,
    CEINMODE,
    CEM,
    CEP,
    CLK,
    C,
    D,
    INMODE,
    MULTSIGNIN,
    OPMODE,
    PCIN,
    RSTA,
    RSTALLCARRYIN,
    RSTALUMODE,
    RSTB,
    RSTC,
    RSTCTRL,
    RSTD,
    RSTINMODE,
    RSTM,
    RSTP);
  output [29:0]ACOUT;
  output [17:0]BCOUT;
  output CARRYCASCOUT;
  output [3:0]CARRYOUT;
  output MULTSIGNOUT;
  output OVERFLOW;
  output PATTERNBDETECT;
  output PATTERNDETECT;
  output [47:0]PCOUT;
  output [47:0]P;
  output UNDERFLOW;
  output [7:0]XOROUT;
  input [29:0]ACIN;
  input [3:0]ALUMODE;
  input [29:0]A;
  input [17:0]BCIN;
  input [17:0]B;
  input CARRYCASCIN;
  input CARRYIN;
  input [2:0]CARRYINSEL;
  input CEA1;
  input CEA2;
  input CEAD;
  input CEALUMODE;
  input CEB1;
  input CEB2;
  input CEC;
  input CECARRYIN;
  input CECTRL;
  input CED;
  input CEINMODE;
  input CEM;
  input CEP;
  input CLK;
  input [47:0]C;
  input [26:0]D;
  input [4:0]INMODE;
  input MULTSIGNIN;
  input [8:0]OPMODE;
  input [47:0]PCIN;
  input RSTA;
  input RSTALLCARRYIN;
  input RSTALUMODE;
  input RSTB;
  input RSTC;
  input RSTCTRL;
  input RSTD;
  input RSTINMODE;
  input RSTM;
  input RSTP;

  wire \ACIN[0] ;
  wire \ACIN[10] ;
  wire \ACIN[11] ;
  wire \ACIN[12] ;
  wire \ACIN[13] ;
  wire \ACIN[14] ;
  wire \ACIN[15] ;
  wire \ACIN[16] ;
  wire \ACIN[17] ;
  wire \ACIN[18] ;
  wire \ACIN[19] ;
  wire \ACIN[1] ;
  wire \ACIN[20] ;
  wire \ACIN[21] ;
  wire \ACIN[22] ;
  wire \ACIN[23] ;
  wire \ACIN[24] ;
  wire \ACIN[25] ;
  wire \ACIN[26] ;
  wire \ACIN[27] ;
  wire \ACIN[28] ;
  wire \ACIN[29] ;
  wire \ACIN[2] ;
  wire \ACIN[3] ;
  wire \ACIN[4] ;
  wire \ACIN[5] ;
  wire \ACIN[6] ;
  wire \ACIN[7] ;
  wire \ACIN[8] ;
  wire \ACIN[9] ;
  wire \ACOUT[0] ;
  wire \ACOUT[10] ;
  wire \ACOUT[11] ;
  wire \ACOUT[12] ;
  wire \ACOUT[13] ;
  wire \ACOUT[14] ;
  wire \ACOUT[15] ;
  wire \ACOUT[16] ;
  wire \ACOUT[17] ;
  wire \ACOUT[18] ;
  wire \ACOUT[19] ;
  wire \ACOUT[1] ;
  wire \ACOUT[20] ;
  wire \ACOUT[21] ;
  wire \ACOUT[22] ;
  wire \ACOUT[23] ;
  wire \ACOUT[24] ;
  wire \ACOUT[25] ;
  wire \ACOUT[26] ;
  wire \ACOUT[27] ;
  wire \ACOUT[28] ;
  wire \ACOUT[29] ;
  wire \ACOUT[2] ;
  wire \ACOUT[3] ;
  wire \ACOUT[4] ;
  wire \ACOUT[5] ;
  wire \ACOUT[6] ;
  wire \ACOUT[7] ;
  wire \ACOUT[8] ;
  wire \ACOUT[9] ;
  wire \ALUMODE[0] ;
  wire \ALUMODE[1] ;
  wire \ALUMODE[2] ;
  wire \ALUMODE[3] ;
  wire \A[0] ;
  wire \A[10] ;
  wire \A[11] ;
  wire \A[12] ;
  wire \A[13] ;
  wire \A[14] ;
  wire \A[15] ;
  wire \A[16] ;
  wire \A[17] ;
  wire \A[18] ;
  wire \A[19] ;
  wire \A[1] ;
  wire \A[20] ;
  wire \A[21] ;
  wire \A[22] ;
  wire \A[23] ;
  wire \A[24] ;
  wire \A[25] ;
  wire \A[26] ;
  wire \A[27] ;
  wire \A[28] ;
  wire \A[29] ;
  wire \A[2] ;
  wire \A[3] ;
  wire \A[4] ;
  wire \A[5] ;
  wire \A[6] ;
  wire \A[7] ;
  wire \A[8] ;
  wire \A[9] ;
  wire \BCIN[0] ;
  wire \BCIN[10] ;
  wire \BCIN[11] ;
  wire \BCIN[12] ;
  wire \BCIN[13] ;
  wire \BCIN[14] ;
  wire \BCIN[15] ;
  wire \BCIN[16] ;
  wire \BCIN[17] ;
  wire \BCIN[1] ;
  wire \BCIN[2] ;
  wire \BCIN[3] ;
  wire \BCIN[4] ;
  wire \BCIN[5] ;
  wire \BCIN[6] ;
  wire \BCIN[7] ;
  wire \BCIN[8] ;
  wire \BCIN[9] ;
  wire \BCOUT[0] ;
  wire \BCOUT[10] ;
  wire \BCOUT[11] ;
  wire \BCOUT[12] ;
  wire \BCOUT[13] ;
  wire \BCOUT[14] ;
  wire \BCOUT[15] ;
  wire \BCOUT[16] ;
  wire \BCOUT[17] ;
  wire \BCOUT[1] ;
  wire \BCOUT[2] ;
  wire \BCOUT[3] ;
  wire \BCOUT[4] ;
  wire \BCOUT[5] ;
  wire \BCOUT[6] ;
  wire \BCOUT[7] ;
  wire \BCOUT[8] ;
  wire \BCOUT[9] ;
  wire \B[0] ;
  wire \B[10] ;
  wire \B[11] ;
  wire \B[12] ;
  wire \B[13] ;
  wire \B[14] ;
  wire \B[15] ;
  wire \B[16] ;
  wire \B[17] ;
  wire \B[1] ;
  wire \B[2] ;
  wire \B[3] ;
  wire \B[4] ;
  wire \B[5] ;
  wire \B[6] ;
  wire \B[7] ;
  wire \B[8] ;
  wire \B[9] ;
  wire CARRYCASCIN;
  wire CARRYCASCOUT;
  wire CARRYIN;
  wire \CARRYINSEL[0] ;
  wire \CARRYINSEL[1] ;
  wire \CARRYINSEL[2] ;
  wire \CARRYOUT[0] ;
  wire \CARRYOUT[1] ;
  wire \CARRYOUT[2] ;
  wire \CARRYOUT[3] ;
  wire CEA1;
  wire CEA2;
  wire CEAD;
  wire CEALUMODE;
  wire CEB1;
  wire CEB2;
  wire CEC;
  wire CECARRYIN;
  wire CECTRL;
  wire CED;
  wire CEINMODE;
  wire CEM;
  wire CEP;
  wire CLK;
  wire \C[0] ;
  wire \C[10] ;
  wire \C[11] ;
  wire \C[12] ;
  wire \C[13] ;
  wire \C[14] ;
  wire \C[15] ;
  wire \C[16] ;
  wire \C[17] ;
  wire \C[18] ;
  wire \C[19] ;
  wire \C[1] ;
  wire \C[20] ;
  wire \C[21] ;
  wire \C[22] ;
  wire \C[23] ;
  wire \C[24] ;
  wire \C[25] ;
  wire \C[26] ;
  wire \C[27] ;
  wire \C[28] ;
  wire \C[29] ;
  wire \C[2] ;
  wire \C[30] ;
  wire \C[31] ;
  wire \C[32] ;
  wire \C[33] ;
  wire \C[34] ;
  wire \C[35] ;
  wire \C[36] ;
  wire \C[37] ;
  wire \C[38] ;
  wire \C[39] ;
  wire \C[3] ;
  wire \C[40] ;
  wire \C[41] ;
  wire \C[42] ;
  wire \C[43] ;
  wire \C[44] ;
  wire \C[45] ;
  wire \C[46] ;
  wire \C[47] ;
  wire \C[4] ;
  wire \C[5] ;
  wire \C[6] ;
  wire \C[7] ;
  wire \C[8] ;
  wire \C[9] ;
  wire \DSP_ALU.ALUMODE10 ;
  wire \DSP_ALU.ALU_OUT<0> ;
  wire \DSP_ALU.ALU_OUT<10> ;
  wire \DSP_ALU.ALU_OUT<11> ;
  wire \DSP_ALU.ALU_OUT<12> ;
  wire \DSP_ALU.ALU_OUT<13> ;
  wire \DSP_ALU.ALU_OUT<14> ;
  wire \DSP_ALU.ALU_OUT<15> ;
  wire \DSP_ALU.ALU_OUT<16> ;
  wire \DSP_ALU.ALU_OUT<17> ;
  wire \DSP_ALU.ALU_OUT<18> ;
  wire \DSP_ALU.ALU_OUT<19> ;
  wire \DSP_ALU.ALU_OUT<1> ;
  wire \DSP_ALU.ALU_OUT<20> ;
  wire \DSP_ALU.ALU_OUT<21> ;
  wire \DSP_ALU.ALU_OUT<22> ;
  wire \DSP_ALU.ALU_OUT<23> ;
  wire \DSP_ALU.ALU_OUT<24> ;
  wire \DSP_ALU.ALU_OUT<25> ;
  wire \DSP_ALU.ALU_OUT<26> ;
  wire \DSP_ALU.ALU_OUT<27> ;
  wire \DSP_ALU.ALU_OUT<28> ;
  wire \DSP_ALU.ALU_OUT<29> ;
  wire \DSP_ALU.ALU_OUT<2> ;
  wire \DSP_ALU.ALU_OUT<30> ;
  wire \DSP_ALU.ALU_OUT<31> ;
  wire \DSP_ALU.ALU_OUT<32> ;
  wire \DSP_ALU.ALU_OUT<33> ;
  wire \DSP_ALU.ALU_OUT<34> ;
  wire \DSP_ALU.ALU_OUT<35> ;
  wire \DSP_ALU.ALU_OUT<36> ;
  wire \DSP_ALU.ALU_OUT<37> ;
  wire \DSP_ALU.ALU_OUT<38> ;
  wire \DSP_ALU.ALU_OUT<39> ;
  wire \DSP_ALU.ALU_OUT<3> ;
  wire \DSP_ALU.ALU_OUT<40> ;
  wire \DSP_ALU.ALU_OUT<41> ;
  wire \DSP_ALU.ALU_OUT<42> ;
  wire \DSP_ALU.ALU_OUT<43> ;
  wire \DSP_ALU.ALU_OUT<44> ;
  wire \DSP_ALU.ALU_OUT<45> ;
  wire \DSP_ALU.ALU_OUT<46> ;
  wire \DSP_ALU.ALU_OUT<47> ;
  wire \DSP_ALU.ALU_OUT<4> ;
  wire \DSP_ALU.ALU_OUT<5> ;
  wire \DSP_ALU.ALU_OUT<6> ;
  wire \DSP_ALU.ALU_OUT<7> ;
  wire \DSP_ALU.ALU_OUT<8> ;
  wire \DSP_ALU.ALU_OUT<9> ;
  wire \DSP_ALU.COUT<0> ;
  wire \DSP_ALU.COUT<1> ;
  wire \DSP_ALU.COUT<2> ;
  wire \DSP_ALU.COUT<3> ;
  wire \DSP_ALU.MULTSIGN_ALU ;
  wire \DSP_ALU.XOR_MX<0> ;
  wire \DSP_ALU.XOR_MX<1> ;
  wire \DSP_ALU.XOR_MX<2> ;
  wire \DSP_ALU.XOR_MX<3> ;
  wire \DSP_ALU.XOR_MX<4> ;
  wire \DSP_ALU.XOR_MX<5> ;
  wire \DSP_ALU.XOR_MX<6> ;
  wire \DSP_ALU.XOR_MX<7> ;
  wire \DSP_A_B_DATA.A1_DATA<0> ;
  wire \DSP_A_B_DATA.A1_DATA<10> ;
  wire \DSP_A_B_DATA.A1_DATA<11> ;
  wire \DSP_A_B_DATA.A1_DATA<12> ;
  wire \DSP_A_B_DATA.A1_DATA<13> ;
  wire \DSP_A_B_DATA.A1_DATA<14> ;
  wire \DSP_A_B_DATA.A1_DATA<15> ;
  wire \DSP_A_B_DATA.A1_DATA<16> ;
  wire \DSP_A_B_DATA.A1_DATA<17> ;
  wire \DSP_A_B_DATA.A1_DATA<18> ;
  wire \DSP_A_B_DATA.A1_DATA<19> ;
  wire \DSP_A_B_DATA.A1_DATA<1> ;
  wire \DSP_A_B_DATA.A1_DATA<20> ;
  wire \DSP_A_B_DATA.A1_DATA<21> ;
  wire \DSP_A_B_DATA.A1_DATA<22> ;
  wire \DSP_A_B_DATA.A1_DATA<23> ;
  wire \DSP_A_B_DATA.A1_DATA<24> ;
  wire \DSP_A_B_DATA.A1_DATA<25> ;
  wire \DSP_A_B_DATA.A1_DATA<26> ;
  wire \DSP_A_B_DATA.A1_DATA<2> ;
  wire \DSP_A_B_DATA.A1_DATA<3> ;
  wire \DSP_A_B_DATA.A1_DATA<4> ;
  wire \DSP_A_B_DATA.A1_DATA<5> ;
  wire \DSP_A_B_DATA.A1_DATA<6> ;
  wire \DSP_A_B_DATA.A1_DATA<7> ;
  wire \DSP_A_B_DATA.A1_DATA<8> ;
  wire \DSP_A_B_DATA.A1_DATA<9> ;
  wire \DSP_A_B_DATA.A2_DATA<0> ;
  wire \DSP_A_B_DATA.A2_DATA<10> ;
  wire \DSP_A_B_DATA.A2_DATA<11> ;
  wire \DSP_A_B_DATA.A2_DATA<12> ;
  wire \DSP_A_B_DATA.A2_DATA<13> ;
  wire \DSP_A_B_DATA.A2_DATA<14> ;
  wire \DSP_A_B_DATA.A2_DATA<15> ;
  wire \DSP_A_B_DATA.A2_DATA<16> ;
  wire \DSP_A_B_DATA.A2_DATA<17> ;
  wire \DSP_A_B_DATA.A2_DATA<18> ;
  wire \DSP_A_B_DATA.A2_DATA<19> ;
  wire \DSP_A_B_DATA.A2_DATA<1> ;
  wire \DSP_A_B_DATA.A2_DATA<20> ;
  wire \DSP_A_B_DATA.A2_DATA<21> ;
  wire \DSP_A_B_DATA.A2_DATA<22> ;
  wire \DSP_A_B_DATA.A2_DATA<23> ;
  wire \DSP_A_B_DATA.A2_DATA<24> ;
  wire \DSP_A_B_DATA.A2_DATA<25> ;
  wire \DSP_A_B_DATA.A2_DATA<26> ;
  wire \DSP_A_B_DATA.A2_DATA<2> ;
  wire \DSP_A_B_DATA.A2_DATA<3> ;
  wire \DSP_A_B_DATA.A2_DATA<4> ;
  wire \DSP_A_B_DATA.A2_DATA<5> ;
  wire \DSP_A_B_DATA.A2_DATA<6> ;
  wire \DSP_A_B_DATA.A2_DATA<7> ;
  wire \DSP_A_B_DATA.A2_DATA<8> ;
  wire \DSP_A_B_DATA.A2_DATA<9> ;
  wire \DSP_A_B_DATA.A_ALU<0> ;
  wire \DSP_A_B_DATA.A_ALU<10> ;
  wire \DSP_A_B_DATA.A_ALU<11> ;
  wire \DSP_A_B_DATA.A_ALU<12> ;
  wire \DSP_A_B_DATA.A_ALU<13> ;
  wire \DSP_A_B_DATA.A_ALU<14> ;
  wire \DSP_A_B_DATA.A_ALU<15> ;
  wire \DSP_A_B_DATA.A_ALU<16> ;
  wire \DSP_A_B_DATA.A_ALU<17> ;
  wire \DSP_A_B_DATA.A_ALU<18> ;
  wire \DSP_A_B_DATA.A_ALU<19> ;
  wire \DSP_A_B_DATA.A_ALU<1> ;
  wire \DSP_A_B_DATA.A_ALU<20> ;
  wire \DSP_A_B_DATA.A_ALU<21> ;
  wire \DSP_A_B_DATA.A_ALU<22> ;
  wire \DSP_A_B_DATA.A_ALU<23> ;
  wire \DSP_A_B_DATA.A_ALU<24> ;
  wire \DSP_A_B_DATA.A_ALU<25> ;
  wire \DSP_A_B_DATA.A_ALU<26> ;
  wire \DSP_A_B_DATA.A_ALU<27> ;
  wire \DSP_A_B_DATA.A_ALU<28> ;
  wire \DSP_A_B_DATA.A_ALU<29> ;
  wire \DSP_A_B_DATA.A_ALU<2> ;
  wire \DSP_A_B_DATA.A_ALU<3> ;
  wire \DSP_A_B_DATA.A_ALU<4> ;
  wire \DSP_A_B_DATA.A_ALU<5> ;
  wire \DSP_A_B_DATA.A_ALU<6> ;
  wire \DSP_A_B_DATA.A_ALU<7> ;
  wire \DSP_A_B_DATA.A_ALU<8> ;
  wire \DSP_A_B_DATA.A_ALU<9> ;
  wire \DSP_A_B_DATA.B1_DATA<0> ;
  wire \DSP_A_B_DATA.B1_DATA<10> ;
  wire \DSP_A_B_DATA.B1_DATA<11> ;
  wire \DSP_A_B_DATA.B1_DATA<12> ;
  wire \DSP_A_B_DATA.B1_DATA<13> ;
  wire \DSP_A_B_DATA.B1_DATA<14> ;
  wire \DSP_A_B_DATA.B1_DATA<15> ;
  wire \DSP_A_B_DATA.B1_DATA<16> ;
  wire \DSP_A_B_DATA.B1_DATA<17> ;
  wire \DSP_A_B_DATA.B1_DATA<1> ;
  wire \DSP_A_B_DATA.B1_DATA<2> ;
  wire \DSP_A_B_DATA.B1_DATA<3> ;
  wire \DSP_A_B_DATA.B1_DATA<4> ;
  wire \DSP_A_B_DATA.B1_DATA<5> ;
  wire \DSP_A_B_DATA.B1_DATA<6> ;
  wire \DSP_A_B_DATA.B1_DATA<7> ;
  wire \DSP_A_B_DATA.B1_DATA<8> ;
  wire \DSP_A_B_DATA.B1_DATA<9> ;
  wire \DSP_A_B_DATA.B2_DATA<0> ;
  wire \DSP_A_B_DATA.B2_DATA<10> ;
  wire \DSP_A_B_DATA.B2_DATA<11> ;
  wire \DSP_A_B_DATA.B2_DATA<12> ;
  wire \DSP_A_B_DATA.B2_DATA<13> ;
  wire \DSP_A_B_DATA.B2_DATA<14> ;
  wire \DSP_A_B_DATA.B2_DATA<15> ;
  wire \DSP_A_B_DATA.B2_DATA<16> ;
  wire \DSP_A_B_DATA.B2_DATA<17> ;
  wire \DSP_A_B_DATA.B2_DATA<1> ;
  wire \DSP_A_B_DATA.B2_DATA<2> ;
  wire \DSP_A_B_DATA.B2_DATA<3> ;
  wire \DSP_A_B_DATA.B2_DATA<4> ;
  wire \DSP_A_B_DATA.B2_DATA<5> ;
  wire \DSP_A_B_DATA.B2_DATA<6> ;
  wire \DSP_A_B_DATA.B2_DATA<7> ;
  wire \DSP_A_B_DATA.B2_DATA<8> ;
  wire \DSP_A_B_DATA.B2_DATA<9> ;
  wire \DSP_A_B_DATA.B_ALU<0> ;
  wire \DSP_A_B_DATA.B_ALU<10> ;
  wire \DSP_A_B_DATA.B_ALU<11> ;
  wire \DSP_A_B_DATA.B_ALU<12> ;
  wire \DSP_A_B_DATA.B_ALU<13> ;
  wire \DSP_A_B_DATA.B_ALU<14> ;
  wire \DSP_A_B_DATA.B_ALU<15> ;
  wire \DSP_A_B_DATA.B_ALU<16> ;
  wire \DSP_A_B_DATA.B_ALU<17> ;
  wire \DSP_A_B_DATA.B_ALU<1> ;
  wire \DSP_A_B_DATA.B_ALU<2> ;
  wire \DSP_A_B_DATA.B_ALU<3> ;
  wire \DSP_A_B_DATA.B_ALU<4> ;
  wire \DSP_A_B_DATA.B_ALU<5> ;
  wire \DSP_A_B_DATA.B_ALU<6> ;
  wire \DSP_A_B_DATA.B_ALU<7> ;
  wire \DSP_A_B_DATA.B_ALU<8> ;
  wire \DSP_A_B_DATA.B_ALU<9> ;
  wire \DSP_C_DATA.C_DATA<0> ;
  wire \DSP_C_DATA.C_DATA<10> ;
  wire \DSP_C_DATA.C_DATA<11> ;
  wire \DSP_C_DATA.C_DATA<12> ;
  wire \DSP_C_DATA.C_DATA<13> ;
  wire \DSP_C_DATA.C_DATA<14> ;
  wire \DSP_C_DATA.C_DATA<15> ;
  wire \DSP_C_DATA.C_DATA<16> ;
  wire \DSP_C_DATA.C_DATA<17> ;
  wire \DSP_C_DATA.C_DATA<18> ;
  wire \DSP_C_DATA.C_DATA<19> ;
  wire \DSP_C_DATA.C_DATA<1> ;
  wire \DSP_C_DATA.C_DATA<20> ;
  wire \DSP_C_DATA.C_DATA<21> ;
  wire \DSP_C_DATA.C_DATA<22> ;
  wire \DSP_C_DATA.C_DATA<23> ;
  wire \DSP_C_DATA.C_DATA<24> ;
  wire \DSP_C_DATA.C_DATA<25> ;
  wire \DSP_C_DATA.C_DATA<26> ;
  wire \DSP_C_DATA.C_DATA<27> ;
  wire \DSP_C_DATA.C_DATA<28> ;
  wire \DSP_C_DATA.C_DATA<29> ;
  wire \DSP_C_DATA.C_DATA<2> ;
  wire \DSP_C_DATA.C_DATA<30> ;
  wire \DSP_C_DATA.C_DATA<31> ;
  wire \DSP_C_DATA.C_DATA<32> ;
  wire \DSP_C_DATA.C_DATA<33> ;
  wire \DSP_C_DATA.C_DATA<34> ;
  wire \DSP_C_DATA.C_DATA<35> ;
  wire \DSP_C_DATA.C_DATA<36> ;
  wire \DSP_C_DATA.C_DATA<37> ;
  wire \DSP_C_DATA.C_DATA<38> ;
  wire \DSP_C_DATA.C_DATA<39> ;
  wire \DSP_C_DATA.C_DATA<3> ;
  wire \DSP_C_DATA.C_DATA<40> ;
  wire \DSP_C_DATA.C_DATA<41> ;
  wire \DSP_C_DATA.C_DATA<42> ;
  wire \DSP_C_DATA.C_DATA<43> ;
  wire \DSP_C_DATA.C_DATA<44> ;
  wire \DSP_C_DATA.C_DATA<45> ;
  wire \DSP_C_DATA.C_DATA<46> ;
  wire \DSP_C_DATA.C_DATA<47> ;
  wire \DSP_C_DATA.C_DATA<4> ;
  wire \DSP_C_DATA.C_DATA<5> ;
  wire \DSP_C_DATA.C_DATA<6> ;
  wire \DSP_C_DATA.C_DATA<7> ;
  wire \DSP_C_DATA.C_DATA<8> ;
  wire \DSP_C_DATA.C_DATA<9> ;
  wire \DSP_MULTIPLIER.AMULT26 ;
  wire \DSP_MULTIPLIER.BMULT17 ;
  wire \DSP_MULTIPLIER.U<0> ;
  wire \DSP_MULTIPLIER.U<10> ;
  wire \DSP_MULTIPLIER.U<11> ;
  wire \DSP_MULTIPLIER.U<12> ;
  wire \DSP_MULTIPLIER.U<13> ;
  wire \DSP_MULTIPLIER.U<14> ;
  wire \DSP_MULTIPLIER.U<15> ;
  wire \DSP_MULTIPLIER.U<16> ;
  wire \DSP_MULTIPLIER.U<17> ;
  wire \DSP_MULTIPLIER.U<18> ;
  wire \DSP_MULTIPLIER.U<19> ;
  wire \DSP_MULTIPLIER.U<1> ;
  wire \DSP_MULTIPLIER.U<20> ;
  wire \DSP_MULTIPLIER.U<21> ;
  wire \DSP_MULTIPLIER.U<22> ;
  wire \DSP_MULTIPLIER.U<23> ;
  wire \DSP_MULTIPLIER.U<24> ;
  wire \DSP_MULTIPLIER.U<25> ;
  wire \DSP_MULTIPLIER.U<26> ;
  wire \DSP_MULTIPLIER.U<27> ;
  wire \DSP_MULTIPLIER.U<28> ;
  wire \DSP_MULTIPLIER.U<29> ;
  wire \DSP_MULTIPLIER.U<2> ;
  wire \DSP_MULTIPLIER.U<30> ;
  wire \DSP_MULTIPLIER.U<31> ;
  wire \DSP_MULTIPLIER.U<32> ;
  wire \DSP_MULTIPLIER.U<33> ;
  wire \DSP_MULTIPLIER.U<34> ;
  wire \DSP_MULTIPLIER.U<35> ;
  wire \DSP_MULTIPLIER.U<36> ;
  wire \DSP_MULTIPLIER.U<37> ;
  wire \DSP_MULTIPLIER.U<38> ;
  wire \DSP_MULTIPLIER.U<39> ;
  wire \DSP_MULTIPLIER.U<3> ;
  wire \DSP_MULTIPLIER.U<40> ;
  wire \DSP_MULTIPLIER.U<41> ;
  wire \DSP_MULTIPLIER.U<42> ;
  wire \DSP_MULTIPLIER.U<43> ;
  wire \DSP_MULTIPLIER.U<44> ;
  wire \DSP_MULTIPLIER.U<4> ;
  wire \DSP_MULTIPLIER.U<5> ;
  wire \DSP_MULTIPLIER.U<6> ;
  wire \DSP_MULTIPLIER.U<7> ;
  wire \DSP_MULTIPLIER.U<8> ;
  wire \DSP_MULTIPLIER.U<9> ;
  wire \DSP_MULTIPLIER.V<0> ;
  wire \DSP_MULTIPLIER.V<10> ;
  wire \DSP_MULTIPLIER.V<11> ;
  wire \DSP_MULTIPLIER.V<12> ;
  wire \DSP_MULTIPLIER.V<13> ;
  wire \DSP_MULTIPLIER.V<14> ;
  wire \DSP_MULTIPLIER.V<15> ;
  wire \DSP_MULTIPLIER.V<16> ;
  wire \DSP_MULTIPLIER.V<17> ;
  wire \DSP_MULTIPLIER.V<18> ;
  wire \DSP_MULTIPLIER.V<19> ;
  wire \DSP_MULTIPLIER.V<1> ;
  wire \DSP_MULTIPLIER.V<20> ;
  wire \DSP_MULTIPLIER.V<21> ;
  wire \DSP_MULTIPLIER.V<22> ;
  wire \DSP_MULTIPLIER.V<23> ;
  wire \DSP_MULTIPLIER.V<24> ;
  wire \DSP_MULTIPLIER.V<25> ;
  wire \DSP_MULTIPLIER.V<26> ;
  wire \DSP_MULTIPLIER.V<27> ;
  wire \DSP_MULTIPLIER.V<28> ;
  wire \DSP_MULTIPLIER.V<29> ;
  wire \DSP_MULTIPLIER.V<2> ;
  wire \DSP_MULTIPLIER.V<30> ;
  wire \DSP_MULTIPLIER.V<31> ;
  wire \DSP_MULTIPLIER.V<32> ;
  wire \DSP_MULTIPLIER.V<33> ;
  wire \DSP_MULTIPLIER.V<34> ;
  wire \DSP_MULTIPLIER.V<35> ;
  wire \DSP_MULTIPLIER.V<36> ;
  wire \DSP_MULTIPLIER.V<37> ;
  wire \DSP_MULTIPLIER.V<38> ;
  wire \DSP_MULTIPLIER.V<39> ;
  wire \DSP_MULTIPLIER.V<3> ;
  wire \DSP_MULTIPLIER.V<40> ;
  wire \DSP_MULTIPLIER.V<41> ;
  wire \DSP_MULTIPLIER.V<42> ;
  wire \DSP_MULTIPLIER.V<43> ;
  wire \DSP_MULTIPLIER.V<44> ;
  wire \DSP_MULTIPLIER.V<4> ;
  wire \DSP_MULTIPLIER.V<5> ;
  wire \DSP_MULTIPLIER.V<6> ;
  wire \DSP_MULTIPLIER.V<7> ;
  wire \DSP_MULTIPLIER.V<8> ;
  wire \DSP_MULTIPLIER.V<9> ;
  wire \DSP_M_DATA.U_DATA<0> ;
  wire \DSP_M_DATA.U_DATA<10> ;
  wire \DSP_M_DATA.U_DATA<11> ;
  wire \DSP_M_DATA.U_DATA<12> ;
  wire \DSP_M_DATA.U_DATA<13> ;
  wire \DSP_M_DATA.U_DATA<14> ;
  wire \DSP_M_DATA.U_DATA<15> ;
  wire \DSP_M_DATA.U_DATA<16> ;
  wire \DSP_M_DATA.U_DATA<17> ;
  wire \DSP_M_DATA.U_DATA<18> ;
  wire \DSP_M_DATA.U_DATA<19> ;
  wire \DSP_M_DATA.U_DATA<1> ;
  wire \DSP_M_DATA.U_DATA<20> ;
  wire \DSP_M_DATA.U_DATA<21> ;
  wire \DSP_M_DATA.U_DATA<22> ;
  wire \DSP_M_DATA.U_DATA<23> ;
  wire \DSP_M_DATA.U_DATA<24> ;
  wire \DSP_M_DATA.U_DATA<25> ;
  wire \DSP_M_DATA.U_DATA<26> ;
  wire \DSP_M_DATA.U_DATA<27> ;
  wire \DSP_M_DATA.U_DATA<28> ;
  wire \DSP_M_DATA.U_DATA<29> ;
  wire \DSP_M_DATA.U_DATA<2> ;
  wire \DSP_M_DATA.U_DATA<30> ;
  wire \DSP_M_DATA.U_DATA<31> ;
  wire \DSP_M_DATA.U_DATA<32> ;
  wire \DSP_M_DATA.U_DATA<33> ;
  wire \DSP_M_DATA.U_DATA<34> ;
  wire \DSP_M_DATA.U_DATA<35> ;
  wire \DSP_M_DATA.U_DATA<36> ;
  wire \DSP_M_DATA.U_DATA<37> ;
  wire \DSP_M_DATA.U_DATA<38> ;
  wire \DSP_M_DATA.U_DATA<39> ;
  wire \DSP_M_DATA.U_DATA<3> ;
  wire \DSP_M_DATA.U_DATA<40> ;
  wire \DSP_M_DATA.U_DATA<41> ;
  wire \DSP_M_DATA.U_DATA<42> ;
  wire \DSP_M_DATA.U_DATA<43> ;
  wire \DSP_M_DATA.U_DATA<44> ;
  wire \DSP_M_DATA.U_DATA<4> ;
  wire \DSP_M_DATA.U_DATA<5> ;
  wire \DSP_M_DATA.U_DATA<6> ;
  wire \DSP_M_DATA.U_DATA<7> ;
  wire \DSP_M_DATA.U_DATA<8> ;
  wire \DSP_M_DATA.U_DATA<9> ;
  wire \DSP_M_DATA.V_DATA<0> ;
  wire \DSP_M_DATA.V_DATA<10> ;
  wire \DSP_M_DATA.V_DATA<11> ;
  wire \DSP_M_DATA.V_DATA<12> ;
  wire \DSP_M_DATA.V_DATA<13> ;
  wire \DSP_M_DATA.V_DATA<14> ;
  wire \DSP_M_DATA.V_DATA<15> ;
  wire \DSP_M_DATA.V_DATA<16> ;
  wire \DSP_M_DATA.V_DATA<17> ;
  wire \DSP_M_DATA.V_DATA<18> ;
  wire \DSP_M_DATA.V_DATA<19> ;
  wire \DSP_M_DATA.V_DATA<1> ;
  wire \DSP_M_DATA.V_DATA<20> ;
  wire \DSP_M_DATA.V_DATA<21> ;
  wire \DSP_M_DATA.V_DATA<22> ;
  wire \DSP_M_DATA.V_DATA<23> ;
  wire \DSP_M_DATA.V_DATA<24> ;
  wire \DSP_M_DATA.V_DATA<25> ;
  wire \DSP_M_DATA.V_DATA<26> ;
  wire \DSP_M_DATA.V_DATA<27> ;
  wire \DSP_M_DATA.V_DATA<28> ;
  wire \DSP_M_DATA.V_DATA<29> ;
  wire \DSP_M_DATA.V_DATA<2> ;
  wire \DSP_M_DATA.V_DATA<30> ;
  wire \DSP_M_DATA.V_DATA<31> ;
  wire \DSP_M_DATA.V_DATA<32> ;
  wire \DSP_M_DATA.V_DATA<33> ;
  wire \DSP_M_DATA.V_DATA<34> ;
  wire \DSP_M_DATA.V_DATA<35> ;
  wire \DSP_M_DATA.V_DATA<36> ;
  wire \DSP_M_DATA.V_DATA<37> ;
  wire \DSP_M_DATA.V_DATA<38> ;
  wire \DSP_M_DATA.V_DATA<39> ;
  wire \DSP_M_DATA.V_DATA<3> ;
  wire \DSP_M_DATA.V_DATA<40> ;
  wire \DSP_M_DATA.V_DATA<41> ;
  wire \DSP_M_DATA.V_DATA<42> ;
  wire \DSP_M_DATA.V_DATA<43> ;
  wire \DSP_M_DATA.V_DATA<44> ;
  wire \DSP_M_DATA.V_DATA<4> ;
  wire \DSP_M_DATA.V_DATA<5> ;
  wire \DSP_M_DATA.V_DATA<6> ;
  wire \DSP_M_DATA.V_DATA<7> ;
  wire \DSP_M_DATA.V_DATA<8> ;
  wire \DSP_M_DATA.V_DATA<9> ;
  wire \DSP_OUTPUT.CCOUT_FB ;
  wire \DSP_OUTPUT.P_FDBK<0> ;
  wire \DSP_OUTPUT.P_FDBK<10> ;
  wire \DSP_OUTPUT.P_FDBK<11> ;
  wire \DSP_OUTPUT.P_FDBK<12> ;
  wire \DSP_OUTPUT.P_FDBK<13> ;
  wire \DSP_OUTPUT.P_FDBK<14> ;
  wire \DSP_OUTPUT.P_FDBK<15> ;
  wire \DSP_OUTPUT.P_FDBK<16> ;
  wire \DSP_OUTPUT.P_FDBK<17> ;
  wire \DSP_OUTPUT.P_FDBK<18> ;
  wire \DSP_OUTPUT.P_FDBK<19> ;
  wire \DSP_OUTPUT.P_FDBK<1> ;
  wire \DSP_OUTPUT.P_FDBK<20> ;
  wire \DSP_OUTPUT.P_FDBK<21> ;
  wire \DSP_OUTPUT.P_FDBK<22> ;
  wire \DSP_OUTPUT.P_FDBK<23> ;
  wire \DSP_OUTPUT.P_FDBK<24> ;
  wire \DSP_OUTPUT.P_FDBK<25> ;
  wire \DSP_OUTPUT.P_FDBK<26> ;
  wire \DSP_OUTPUT.P_FDBK<27> ;
  wire \DSP_OUTPUT.P_FDBK<28> ;
  wire \DSP_OUTPUT.P_FDBK<29> ;
  wire \DSP_OUTPUT.P_FDBK<2> ;
  wire \DSP_OUTPUT.P_FDBK<30> ;
  wire \DSP_OUTPUT.P_FDBK<31> ;
  wire \DSP_OUTPUT.P_FDBK<32> ;
  wire \DSP_OUTPUT.P_FDBK<33> ;
  wire \DSP_OUTPUT.P_FDBK<34> ;
  wire \DSP_OUTPUT.P_FDBK<35> ;
  wire \DSP_OUTPUT.P_FDBK<36> ;
  wire \DSP_OUTPUT.P_FDBK<37> ;
  wire \DSP_OUTPUT.P_FDBK<38> ;
  wire \DSP_OUTPUT.P_FDBK<39> ;
  wire \DSP_OUTPUT.P_FDBK<3> ;
  wire \DSP_OUTPUT.P_FDBK<40> ;
  wire \DSP_OUTPUT.P_FDBK<41> ;
  wire \DSP_OUTPUT.P_FDBK<42> ;
  wire \DSP_OUTPUT.P_FDBK<43> ;
  wire \DSP_OUTPUT.P_FDBK<44> ;
  wire \DSP_OUTPUT.P_FDBK<45> ;
  wire \DSP_OUTPUT.P_FDBK<46> ;
  wire \DSP_OUTPUT.P_FDBK<47> ;
  wire \DSP_OUTPUT.P_FDBK<4> ;
  wire \DSP_OUTPUT.P_FDBK<5> ;
  wire \DSP_OUTPUT.P_FDBK<6> ;
  wire \DSP_OUTPUT.P_FDBK<7> ;
  wire \DSP_OUTPUT.P_FDBK<8> ;
  wire \DSP_OUTPUT.P_FDBK<9> ;
  wire \DSP_OUTPUT.P_FDBK_47 ;
  wire \DSP_PREADD.AD<0> ;
  wire \DSP_PREADD.AD<10> ;
  wire \DSP_PREADD.AD<11> ;
  wire \DSP_PREADD.AD<12> ;
  wire \DSP_PREADD.AD<13> ;
  wire \DSP_PREADD.AD<14> ;
  wire \DSP_PREADD.AD<15> ;
  wire \DSP_PREADD.AD<16> ;
  wire \DSP_PREADD.AD<17> ;
  wire \DSP_PREADD.AD<18> ;
  wire \DSP_PREADD.AD<19> ;
  wire \DSP_PREADD.AD<1> ;
  wire \DSP_PREADD.AD<20> ;
  wire \DSP_PREADD.AD<21> ;
  wire \DSP_PREADD.AD<22> ;
  wire \DSP_PREADD.AD<23> ;
  wire \DSP_PREADD.AD<24> ;
  wire \DSP_PREADD.AD<25> ;
  wire \DSP_PREADD.AD<26> ;
  wire \DSP_PREADD.AD<2> ;
  wire \DSP_PREADD.AD<3> ;
  wire \DSP_PREADD.AD<4> ;
  wire \DSP_PREADD.AD<5> ;
  wire \DSP_PREADD.AD<6> ;
  wire \DSP_PREADD.AD<7> ;
  wire \DSP_PREADD.AD<8> ;
  wire \DSP_PREADD.AD<9> ;
  wire \DSP_PREADD_DATA.A2A1<0> ;
  wire \DSP_PREADD_DATA.A2A1<10> ;
  wire \DSP_PREADD_DATA.A2A1<11> ;
  wire \DSP_PREADD_DATA.A2A1<12> ;
  wire \DSP_PREADD_DATA.A2A1<13> ;
  wire \DSP_PREADD_DATA.A2A1<14> ;
  wire \DSP_PREADD_DATA.A2A1<15> ;
  wire \DSP_PREADD_DATA.A2A1<16> ;
  wire \DSP_PREADD_DATA.A2A1<17> ;
  wire \DSP_PREADD_DATA.A2A1<18> ;
  wire \DSP_PREADD_DATA.A2A1<19> ;
  wire \DSP_PREADD_DATA.A2A1<1> ;
  wire \DSP_PREADD_DATA.A2A1<20> ;
  wire \DSP_PREADD_DATA.A2A1<21> ;
  wire \DSP_PREADD_DATA.A2A1<22> ;
  wire \DSP_PREADD_DATA.A2A1<23> ;
  wire \DSP_PREADD_DATA.A2A1<24> ;
  wire \DSP_PREADD_DATA.A2A1<25> ;
  wire \DSP_PREADD_DATA.A2A1<26> ;
  wire \DSP_PREADD_DATA.A2A1<2> ;
  wire \DSP_PREADD_DATA.A2A1<3> ;
  wire \DSP_PREADD_DATA.A2A1<4> ;
  wire \DSP_PREADD_DATA.A2A1<5> ;
  wire \DSP_PREADD_DATA.A2A1<6> ;
  wire \DSP_PREADD_DATA.A2A1<7> ;
  wire \DSP_PREADD_DATA.A2A1<8> ;
  wire \DSP_PREADD_DATA.A2A1<9> ;
  wire \DSP_PREADD_DATA.ADDSUB ;
  wire \DSP_PREADD_DATA.AD_DATA<0> ;
  wire \DSP_PREADD_DATA.AD_DATA<10> ;
  wire \DSP_PREADD_DATA.AD_DATA<11> ;
  wire \DSP_PREADD_DATA.AD_DATA<12> ;
  wire \DSP_PREADD_DATA.AD_DATA<13> ;
  wire \DSP_PREADD_DATA.AD_DATA<14> ;
  wire \DSP_PREADD_DATA.AD_DATA<15> ;
  wire \DSP_PREADD_DATA.AD_DATA<16> ;
  wire \DSP_PREADD_DATA.AD_DATA<17> ;
  wire \DSP_PREADD_DATA.AD_DATA<18> ;
  wire \DSP_PREADD_DATA.AD_DATA<19> ;
  wire \DSP_PREADD_DATA.AD_DATA<1> ;
  wire \DSP_PREADD_DATA.AD_DATA<20> ;
  wire \DSP_PREADD_DATA.AD_DATA<21> ;
  wire \DSP_PREADD_DATA.AD_DATA<22> ;
  wire \DSP_PREADD_DATA.AD_DATA<23> ;
  wire \DSP_PREADD_DATA.AD_DATA<24> ;
  wire \DSP_PREADD_DATA.AD_DATA<25> ;
  wire \DSP_PREADD_DATA.AD_DATA<26> ;
  wire \DSP_PREADD_DATA.AD_DATA<2> ;
  wire \DSP_PREADD_DATA.AD_DATA<3> ;
  wire \DSP_PREADD_DATA.AD_DATA<4> ;
  wire \DSP_PREADD_DATA.AD_DATA<5> ;
  wire \DSP_PREADD_DATA.AD_DATA<6> ;
  wire \DSP_PREADD_DATA.AD_DATA<7> ;
  wire \DSP_PREADD_DATA.AD_DATA<8> ;
  wire \DSP_PREADD_DATA.AD_DATA<9> ;
  wire \DSP_PREADD_DATA.B2B1<0> ;
  wire \DSP_PREADD_DATA.B2B1<10> ;
  wire \DSP_PREADD_DATA.B2B1<11> ;
  wire \DSP_PREADD_DATA.B2B1<12> ;
  wire \DSP_PREADD_DATA.B2B1<13> ;
  wire \DSP_PREADD_DATA.B2B1<14> ;
  wire \DSP_PREADD_DATA.B2B1<15> ;
  wire \DSP_PREADD_DATA.B2B1<16> ;
  wire \DSP_PREADD_DATA.B2B1<17> ;
  wire \DSP_PREADD_DATA.B2B1<1> ;
  wire \DSP_PREADD_DATA.B2B1<2> ;
  wire \DSP_PREADD_DATA.B2B1<3> ;
  wire \DSP_PREADD_DATA.B2B1<4> ;
  wire \DSP_PREADD_DATA.B2B1<5> ;
  wire \DSP_PREADD_DATA.B2B1<6> ;
  wire \DSP_PREADD_DATA.B2B1<7> ;
  wire \DSP_PREADD_DATA.B2B1<8> ;
  wire \DSP_PREADD_DATA.B2B1<9> ;
  wire \DSP_PREADD_DATA.D_DATA<0> ;
  wire \DSP_PREADD_DATA.D_DATA<10> ;
  wire \DSP_PREADD_DATA.D_DATA<11> ;
  wire \DSP_PREADD_DATA.D_DATA<12> ;
  wire \DSP_PREADD_DATA.D_DATA<13> ;
  wire \DSP_PREADD_DATA.D_DATA<14> ;
  wire \DSP_PREADD_DATA.D_DATA<15> ;
  wire \DSP_PREADD_DATA.D_DATA<16> ;
  wire \DSP_PREADD_DATA.D_DATA<17> ;
  wire \DSP_PREADD_DATA.D_DATA<18> ;
  wire \DSP_PREADD_DATA.D_DATA<19> ;
  wire \DSP_PREADD_DATA.D_DATA<1> ;
  wire \DSP_PREADD_DATA.D_DATA<20> ;
  wire \DSP_PREADD_DATA.D_DATA<21> ;
  wire \DSP_PREADD_DATA.D_DATA<22> ;
  wire \DSP_PREADD_DATA.D_DATA<23> ;
  wire \DSP_PREADD_DATA.D_DATA<24> ;
  wire \DSP_PREADD_DATA.D_DATA<25> ;
  wire \DSP_PREADD_DATA.D_DATA<26> ;
  wire \DSP_PREADD_DATA.D_DATA<2> ;
  wire \DSP_PREADD_DATA.D_DATA<3> ;
  wire \DSP_PREADD_DATA.D_DATA<4> ;
  wire \DSP_PREADD_DATA.D_DATA<5> ;
  wire \DSP_PREADD_DATA.D_DATA<6> ;
  wire \DSP_PREADD_DATA.D_DATA<7> ;
  wire \DSP_PREADD_DATA.D_DATA<8> ;
  wire \DSP_PREADD_DATA.D_DATA<9> ;
  wire \DSP_PREADD_DATA.INMODE_2 ;
  wire \DSP_PREADD_DATA.PREADD_AB<0> ;
  wire \DSP_PREADD_DATA.PREADD_AB<10> ;
  wire \DSP_PREADD_DATA.PREADD_AB<11> ;
  wire \DSP_PREADD_DATA.PREADD_AB<12> ;
  wire \DSP_PREADD_DATA.PREADD_AB<13> ;
  wire \DSP_PREADD_DATA.PREADD_AB<14> ;
  wire \DSP_PREADD_DATA.PREADD_AB<15> ;
  wire \DSP_PREADD_DATA.PREADD_AB<16> ;
  wire \DSP_PREADD_DATA.PREADD_AB<17> ;
  wire \DSP_PREADD_DATA.PREADD_AB<18> ;
  wire \DSP_PREADD_DATA.PREADD_AB<19> ;
  wire \DSP_PREADD_DATA.PREADD_AB<1> ;
  wire \DSP_PREADD_DATA.PREADD_AB<20> ;
  wire \DSP_PREADD_DATA.PREADD_AB<21> ;
  wire \DSP_PREADD_DATA.PREADD_AB<22> ;
  wire \DSP_PREADD_DATA.PREADD_AB<23> ;
  wire \DSP_PREADD_DATA.PREADD_AB<24> ;
  wire \DSP_PREADD_DATA.PREADD_AB<25> ;
  wire \DSP_PREADD_DATA.PREADD_AB<26> ;
  wire \DSP_PREADD_DATA.PREADD_AB<2> ;
  wire \DSP_PREADD_DATA.PREADD_AB<3> ;
  wire \DSP_PREADD_DATA.PREADD_AB<4> ;
  wire \DSP_PREADD_DATA.PREADD_AB<5> ;
  wire \DSP_PREADD_DATA.PREADD_AB<6> ;
  wire \DSP_PREADD_DATA.PREADD_AB<7> ;
  wire \DSP_PREADD_DATA.PREADD_AB<8> ;
  wire \DSP_PREADD_DATA.PREADD_AB<9> ;
  wire \D[0] ;
  wire \D[10] ;
  wire \D[11] ;
  wire \D[12] ;
  wire \D[13] ;
  wire \D[14] ;
  wire \D[15] ;
  wire \D[16] ;
  wire \D[17] ;
  wire \D[18] ;
  wire \D[19] ;
  wire \D[1] ;
  wire \D[20] ;
  wire \D[21] ;
  wire \D[22] ;
  wire \D[23] ;
  wire \D[24] ;
  wire \D[25] ;
  wire \D[26] ;
  wire \D[2] ;
  wire \D[3] ;
  wire \D[4] ;
  wire \D[5] ;
  wire \D[6] ;
  wire \D[7] ;
  wire \D[8] ;
  wire \D[9] ;
  wire \INMODE[0] ;
  wire \INMODE[1] ;
  wire \INMODE[2] ;
  wire \INMODE[3] ;
  wire \INMODE[4] ;
  wire MULTSIGNIN;
  wire MULTSIGNOUT;
  wire \OPMODE[0] ;
  wire \OPMODE[1] ;
  wire \OPMODE[2] ;
  wire \OPMODE[3] ;
  wire \OPMODE[4] ;
  wire \OPMODE[5] ;
  wire \OPMODE[6] ;
  wire \OPMODE[7] ;
  wire \OPMODE[8] ;
  wire OVERFLOW;
  wire PATTERNBDETECT;
  wire PATTERNDETECT;
  wire \PCIN[0] ;
  wire \PCIN[10] ;
  wire \PCIN[11] ;
  wire \PCIN[12] ;
  wire \PCIN[13] ;
  wire \PCIN[14] ;
  wire \PCIN[15] ;
  wire \PCIN[16] ;
  wire \PCIN[17] ;
  wire \PCIN[18] ;
  wire \PCIN[19] ;
  wire \PCIN[1] ;
  wire \PCIN[20] ;
  wire \PCIN[21] ;
  wire \PCIN[22] ;
  wire \PCIN[23] ;
  wire \PCIN[24] ;
  wire \PCIN[25] ;
  wire \PCIN[26] ;
  wire \PCIN[27] ;
  wire \PCIN[28] ;
  wire \PCIN[29] ;
  wire \PCIN[2] ;
  wire \PCIN[30] ;
  wire \PCIN[31] ;
  wire \PCIN[32] ;
  wire \PCIN[33] ;
  wire \PCIN[34] ;
  wire \PCIN[35] ;
  wire \PCIN[36] ;
  wire \PCIN[37] ;
  wire \PCIN[38] ;
  wire \PCIN[39] ;
  wire \PCIN[3] ;
  wire \PCIN[40] ;
  wire \PCIN[41] ;
  wire \PCIN[42] ;
  wire \PCIN[43] ;
  wire \PCIN[44] ;
  wire \PCIN[45] ;
  wire \PCIN[46] ;
  wire \PCIN[47] ;
  wire \PCIN[4] ;
  wire \PCIN[5] ;
  wire \PCIN[6] ;
  wire \PCIN[7] ;
  wire \PCIN[8] ;
  wire \PCIN[9] ;
  wire \PCOUT[0] ;
  wire \PCOUT[10] ;
  wire \PCOUT[11] ;
  wire \PCOUT[12] ;
  wire \PCOUT[13] ;
  wire \PCOUT[14] ;
  wire \PCOUT[15] ;
  wire \PCOUT[16] ;
  wire \PCOUT[17] ;
  wire \PCOUT[18] ;
  wire \PCOUT[19] ;
  wire \PCOUT[1] ;
  wire \PCOUT[20] ;
  wire \PCOUT[21] ;
  wire \PCOUT[22] ;
  wire \PCOUT[23] ;
  wire \PCOUT[24] ;
  wire \PCOUT[25] ;
  wire \PCOUT[26] ;
  wire \PCOUT[27] ;
  wire \PCOUT[28] ;
  wire \PCOUT[29] ;
  wire \PCOUT[2] ;
  wire \PCOUT[30] ;
  wire \PCOUT[31] ;
  wire \PCOUT[32] ;
  wire \PCOUT[33] ;
  wire \PCOUT[34] ;
  wire \PCOUT[35] ;
  wire \PCOUT[36] ;
  wire \PCOUT[37] ;
  wire \PCOUT[38] ;
  wire \PCOUT[39] ;
  wire \PCOUT[3] ;
  wire \PCOUT[40] ;
  wire \PCOUT[41] ;
  wire \PCOUT[42] ;
  wire \PCOUT[43] ;
  wire \PCOUT[44] ;
  wire \PCOUT[45] ;
  wire \PCOUT[46] ;
  wire \PCOUT[47] ;
  wire \PCOUT[4] ;
  wire \PCOUT[5] ;
  wire \PCOUT[6] ;
  wire \PCOUT[7] ;
  wire \PCOUT[8] ;
  wire \PCOUT[9] ;
  wire \P[0] ;
  wire \P[10] ;
  wire \P[11] ;
  wire \P[12] ;
  wire \P[13] ;
  wire \P[14] ;
  wire \P[15] ;
  wire \P[16] ;
  wire \P[17] ;
  wire \P[18] ;
  wire \P[19] ;
  wire \P[1] ;
  wire \P[20] ;
  wire \P[21] ;
  wire \P[22] ;
  wire \P[23] ;
  wire \P[24] ;
  wire \P[25] ;
  wire \P[26] ;
  wire \P[27] ;
  wire \P[28] ;
  wire \P[29] ;
  wire \P[2] ;
  wire \P[30] ;
  wire \P[31] ;
  wire \P[32] ;
  wire \P[33] ;
  wire \P[34] ;
  wire \P[35] ;
  wire \P[36] ;
  wire \P[37] ;
  wire \P[38] ;
  wire \P[39] ;
  wire \P[3] ;
  wire \P[40] ;
  wire \P[41] ;
  wire \P[42] ;
  wire \P[43] ;
  wire \P[44] ;
  wire \P[45] ;
  wire \P[46] ;
  wire \P[47] ;
  wire \P[4] ;
  wire \P[5] ;
  wire \P[6] ;
  wire \P[7] ;
  wire \P[8] ;
  wire \P[9] ;
  wire RSTA;
  wire RSTALLCARRYIN;
  wire RSTALUMODE;
  wire RSTB;
  wire RSTC;
  wire RSTCTRL;
  wire RSTD;
  wire RSTINMODE;
  wire RSTM;
  wire RSTP;
  wire UNDERFLOW;
  wire \XOROUT[0] ;
  wire \XOROUT[1] ;
  wire \XOROUT[2] ;
  wire \XOROUT[3] ;
  wire \XOROUT[4] ;
  wire \XOROUT[5] ;
  wire \XOROUT[6] ;
  wire \XOROUT[7] ;

  assign \ACIN[0]  = ACIN[0];
  assign \ACIN[10]  = ACIN[10];
  assign \ACIN[11]  = ACIN[11];
  assign \ACIN[12]  = ACIN[12];
  assign \ACIN[13]  = ACIN[13];
  assign \ACIN[14]  = ACIN[14];
  assign \ACIN[15]  = ACIN[15];
  assign \ACIN[16]  = ACIN[16];
  assign \ACIN[17]  = ACIN[17];
  assign \ACIN[18]  = ACIN[18];
  assign \ACIN[19]  = ACIN[19];
  assign \ACIN[1]  = ACIN[1];
  assign \ACIN[20]  = ACIN[20];
  assign \ACIN[21]  = ACIN[21];
  assign \ACIN[22]  = ACIN[22];
  assign \ACIN[23]  = ACIN[23];
  assign \ACIN[24]  = ACIN[24];
  assign \ACIN[25]  = ACIN[25];
  assign \ACIN[26]  = ACIN[26];
  assign \ACIN[27]  = ACIN[27];
  assign \ACIN[28]  = ACIN[28];
  assign \ACIN[29]  = ACIN[29];
  assign \ACIN[2]  = ACIN[2];
  assign \ACIN[3]  = ACIN[3];
  assign \ACIN[4]  = ACIN[4];
  assign \ACIN[5]  = ACIN[5];
  assign \ACIN[6]  = ACIN[6];
  assign \ACIN[7]  = ACIN[7];
  assign \ACIN[8]  = ACIN[8];
  assign \ACIN[9]  = ACIN[9];
  assign ACOUT[29] = \ACOUT[29] ;
  assign ACOUT[28] = \ACOUT[28] ;
  assign ACOUT[27] = \ACOUT[27] ;
  assign ACOUT[26] = \ACOUT[26] ;
  assign ACOUT[25] = \ACOUT[25] ;
  assign ACOUT[24] = \ACOUT[24] ;
  assign ACOUT[23] = \ACOUT[23] ;
  assign ACOUT[22] = \ACOUT[22] ;
  assign ACOUT[21] = \ACOUT[21] ;
  assign ACOUT[20] = \ACOUT[20] ;
  assign ACOUT[19] = \ACOUT[19] ;
  assign ACOUT[18] = \ACOUT[18] ;
  assign ACOUT[17] = \ACOUT[17] ;
  assign ACOUT[16] = \ACOUT[16] ;
  assign ACOUT[15] = \ACOUT[15] ;
  assign ACOUT[14] = \ACOUT[14] ;
  assign ACOUT[13] = \ACOUT[13] ;
  assign ACOUT[12] = \ACOUT[12] ;
  assign ACOUT[11] = \ACOUT[11] ;
  assign ACOUT[10] = \ACOUT[10] ;
  assign ACOUT[9] = \ACOUT[9] ;
  assign ACOUT[8] = \ACOUT[8] ;
  assign ACOUT[7] = \ACOUT[7] ;
  assign ACOUT[6] = \ACOUT[6] ;
  assign ACOUT[5] = \ACOUT[5] ;
  assign ACOUT[4] = \ACOUT[4] ;
  assign ACOUT[3] = \ACOUT[3] ;
  assign ACOUT[2] = \ACOUT[2] ;
  assign ACOUT[1] = \ACOUT[1] ;
  assign ACOUT[0] = \ACOUT[0] ;
  assign \ALUMODE[0]  = ALUMODE[0];
  assign \ALUMODE[1]  = ALUMODE[1];
  assign \ALUMODE[2]  = ALUMODE[2];
  assign \ALUMODE[3]  = ALUMODE[3];
  assign \A[0]  = A[0];
  assign \A[10]  = A[10];
  assign \A[11]  = A[11];
  assign \A[12]  = A[12];
  assign \A[13]  = A[13];
  assign \A[14]  = A[14];
  assign \A[15]  = A[15];
  assign \A[16]  = A[16];
  assign \A[17]  = A[17];
  assign \A[18]  = A[18];
  assign \A[19]  = A[19];
  assign \A[1]  = A[1];
  assign \A[20]  = A[20];
  assign \A[21]  = A[21];
  assign \A[22]  = A[22];
  assign \A[23]  = A[23];
  assign \A[24]  = A[24];
  assign \A[25]  = A[25];
  assign \A[26]  = A[26];
  assign \A[27]  = A[27];
  assign \A[28]  = A[28];
  assign \A[29]  = A[29];
  assign \A[2]  = A[2];
  assign \A[3]  = A[3];
  assign \A[4]  = A[4];
  assign \A[5]  = A[5];
  assign \A[6]  = A[6];
  assign \A[7]  = A[7];
  assign \A[8]  = A[8];
  assign \A[9]  = A[9];
  assign \BCIN[0]  = BCIN[0];
  assign \BCIN[10]  = BCIN[10];
  assign \BCIN[11]  = BCIN[11];
  assign \BCIN[12]  = BCIN[12];
  assign \BCIN[13]  = BCIN[13];
  assign \BCIN[14]  = BCIN[14];
  assign \BCIN[15]  = BCIN[15];
  assign \BCIN[16]  = BCIN[16];
  assign \BCIN[17]  = BCIN[17];
  assign \BCIN[1]  = BCIN[1];
  assign \BCIN[2]  = BCIN[2];
  assign \BCIN[3]  = BCIN[3];
  assign \BCIN[4]  = BCIN[4];
  assign \BCIN[5]  = BCIN[5];
  assign \BCIN[6]  = BCIN[6];
  assign \BCIN[7]  = BCIN[7];
  assign \BCIN[8]  = BCIN[8];
  assign \BCIN[9]  = BCIN[9];
  assign BCOUT[17] = \BCOUT[17] ;
  assign BCOUT[16] = \BCOUT[16] ;
  assign BCOUT[15] = \BCOUT[15] ;
  assign BCOUT[14] = \BCOUT[14] ;
  assign BCOUT[13] = \BCOUT[13] ;
  assign BCOUT[12] = \BCOUT[12] ;
  assign BCOUT[11] = \BCOUT[11] ;
  assign BCOUT[10] = \BCOUT[10] ;
  assign BCOUT[9] = \BCOUT[9] ;
  assign BCOUT[8] = \BCOUT[8] ;
  assign BCOUT[7] = \BCOUT[7] ;
  assign BCOUT[6] = \BCOUT[6] ;
  assign BCOUT[5] = \BCOUT[5] ;
  assign BCOUT[4] = \BCOUT[4] ;
  assign BCOUT[3] = \BCOUT[3] ;
  assign BCOUT[2] = \BCOUT[2] ;
  assign BCOUT[1] = \BCOUT[1] ;
  assign BCOUT[0] = \BCOUT[0] ;
  assign \B[0]  = B[0];
  assign \B[10]  = B[10];
  assign \B[11]  = B[11];
  assign \B[12]  = B[12];
  assign \B[13]  = B[13];
  assign \B[14]  = B[14];
  assign \B[15]  = B[15];
  assign \B[16]  = B[16];
  assign \B[17]  = B[17];
  assign \B[1]  = B[1];
  assign \B[2]  = B[2];
  assign \B[3]  = B[3];
  assign \B[4]  = B[4];
  assign \B[5]  = B[5];
  assign \B[6]  = B[6];
  assign \B[7]  = B[7];
  assign \B[8]  = B[8];
  assign \B[9]  = B[9];
  assign \CARRYINSEL[0]  = CARRYINSEL[0];
  assign \CARRYINSEL[1]  = CARRYINSEL[1];
  assign \CARRYINSEL[2]  = CARRYINSEL[2];
  assign CARRYOUT[3] = \CARRYOUT[3] ;
  assign CARRYOUT[2] = \CARRYOUT[2] ;
  assign CARRYOUT[1] = \CARRYOUT[1] ;
  assign CARRYOUT[0] = \CARRYOUT[0] ;
  assign \C[0]  = C[0];
  assign \C[10]  = C[10];
  assign \C[11]  = C[11];
  assign \C[12]  = C[12];
  assign \C[13]  = C[13];
  assign \C[14]  = C[14];
  assign \C[15]  = C[15];
  assign \C[16]  = C[16];
  assign \C[17]  = C[17];
  assign \C[18]  = C[18];
  assign \C[19]  = C[19];
  assign \C[1]  = C[1];
  assign \C[20]  = C[20];
  assign \C[21]  = C[21];
  assign \C[22]  = C[22];
  assign \C[23]  = C[23];
  assign \C[24]  = C[24];
  assign \C[25]  = C[25];
  assign \C[26]  = C[26];
  assign \C[27]  = C[27];
  assign \C[28]  = C[28];
  assign \C[29]  = C[29];
  assign \C[2]  = C[2];
  assign \C[30]  = C[30];
  assign \C[31]  = C[31];
  assign \C[32]  = C[32];
  assign \C[33]  = C[33];
  assign \C[34]  = C[34];
  assign \C[35]  = C[35];
  assign \C[36]  = C[36];
  assign \C[37]  = C[37];
  assign \C[38]  = C[38];
  assign \C[39]  = C[39];
  assign \C[3]  = C[3];
  assign \C[40]  = C[40];
  assign \C[41]  = C[41];
  assign \C[42]  = C[42];
  assign \C[43]  = C[43];
  assign \C[44]  = C[44];
  assign \C[45]  = C[45];
  assign \C[46]  = C[46];
  assign \C[47]  = C[47];
  assign \C[4]  = C[4];
  assign \C[5]  = C[5];
  assign \C[6]  = C[6];
  assign \C[7]  = C[7];
  assign \C[8]  = C[8];
  assign \C[9]  = C[9];
  assign \D[0]  = D[0];
  assign \D[10]  = D[10];
  assign \D[11]  = D[11];
  assign \D[12]  = D[12];
  assign \D[13]  = D[13];
  assign \D[14]  = D[14];
  assign \D[15]  = D[15];
  assign \D[16]  = D[16];
  assign \D[17]  = D[17];
  assign \D[18]  = D[18];
  assign \D[19]  = D[19];
  assign \D[1]  = D[1];
  assign \D[20]  = D[20];
  assign \D[21]  = D[21];
  assign \D[22]  = D[22];
  assign \D[23]  = D[23];
  assign \D[24]  = D[24];
  assign \D[25]  = D[25];
  assign \D[26]  = D[26];
  assign \D[2]  = D[2];
  assign \D[3]  = D[3];
  assign \D[4]  = D[4];
  assign \D[5]  = D[5];
  assign \D[6]  = D[6];
  assign \D[7]  = D[7];
  assign \D[8]  = D[8];
  assign \D[9]  = D[9];
  assign \INMODE[0]  = INMODE[0];
  assign \INMODE[1]  = INMODE[1];
  assign \INMODE[2]  = INMODE[2];
  assign \INMODE[3]  = INMODE[3];
  assign \INMODE[4]  = INMODE[4];
  assign \OPMODE[0]  = OPMODE[0];
  assign \OPMODE[1]  = OPMODE[1];
  assign \OPMODE[2]  = OPMODE[2];
  assign \OPMODE[3]  = OPMODE[3];
  assign \OPMODE[4]  = OPMODE[4];
  assign \OPMODE[5]  = OPMODE[5];
  assign \OPMODE[6]  = OPMODE[6];
  assign \OPMODE[7]  = OPMODE[7];
  assign \OPMODE[8]  = OPMODE[8];
  assign P[47] = \P[47] ;
  assign P[46] = \P[46] ;
  assign P[45] = \P[45] ;
  assign P[44] = \P[44] ;
  assign P[43] = \P[43] ;
  assign P[42] = \P[42] ;
  assign P[41] = \P[41] ;
  assign P[40] = \P[40] ;
  assign P[39] = \P[39] ;
  assign P[38] = \P[38] ;
  assign P[37] = \P[37] ;
  assign P[36] = \P[36] ;
  assign P[35] = \P[35] ;
  assign P[34] = \P[34] ;
  assign P[33] = \P[33] ;
  assign P[32] = \P[32] ;
  assign P[31] = \P[31] ;
  assign P[30] = \P[30] ;
  assign P[29] = \P[29] ;
  assign P[28] = \P[28] ;
  assign P[27] = \P[27] ;
  assign P[26] = \P[26] ;
  assign P[25] = \P[25] ;
  assign P[24] = \P[24] ;
  assign P[23] = \P[23] ;
  assign P[22] = \P[22] ;
  assign P[21] = \P[21] ;
  assign P[20] = \P[20] ;
  assign P[19] = \P[19] ;
  assign P[18] = \P[18] ;
  assign P[17] = \P[17] ;
  assign P[16] = \P[16] ;
  assign P[15] = \P[15] ;
  assign P[14] = \P[14] ;
  assign P[13] = \P[13] ;
  assign P[12] = \P[12] ;
  assign P[11] = \P[11] ;
  assign P[10] = \P[10] ;
  assign P[9] = \P[9] ;
  assign P[8] = \P[8] ;
  assign P[7] = \P[7] ;
  assign P[6] = \P[6] ;
  assign P[5] = \P[5] ;
  assign P[4] = \P[4] ;
  assign P[3] = \P[3] ;
  assign P[2] = \P[2] ;
  assign P[1] = \P[1] ;
  assign P[0] = \P[0] ;
  assign \PCIN[0]  = PCIN[0];
  assign \PCIN[10]  = PCIN[10];
  assign \PCIN[11]  = PCIN[11];
  assign \PCIN[12]  = PCIN[12];
  assign \PCIN[13]  = PCIN[13];
  assign \PCIN[14]  = PCIN[14];
  assign \PCIN[15]  = PCIN[15];
  assign \PCIN[16]  = PCIN[16];
  assign \PCIN[17]  = PCIN[17];
  assign \PCIN[18]  = PCIN[18];
  assign \PCIN[19]  = PCIN[19];
  assign \PCIN[1]  = PCIN[1];
  assign \PCIN[20]  = PCIN[20];
  assign \PCIN[21]  = PCIN[21];
  assign \PCIN[22]  = PCIN[22];
  assign \PCIN[23]  = PCIN[23];
  assign \PCIN[24]  = PCIN[24];
  assign \PCIN[25]  = PCIN[25];
  assign \PCIN[26]  = PCIN[26];
  assign \PCIN[27]  = PCIN[27];
  assign \PCIN[28]  = PCIN[28];
  assign \PCIN[29]  = PCIN[29];
  assign \PCIN[2]  = PCIN[2];
  assign \PCIN[30]  = PCIN[30];
  assign \PCIN[31]  = PCIN[31];
  assign \PCIN[32]  = PCIN[32];
  assign \PCIN[33]  = PCIN[33];
  assign \PCIN[34]  = PCIN[34];
  assign \PCIN[35]  = PCIN[35];
  assign \PCIN[36]  = PCIN[36];
  assign \PCIN[37]  = PCIN[37];
  assign \PCIN[38]  = PCIN[38];
  assign \PCIN[39]  = PCIN[39];
  assign \PCIN[3]  = PCIN[3];
  assign \PCIN[40]  = PCIN[40];
  assign \PCIN[41]  = PCIN[41];
  assign \PCIN[42]  = PCIN[42];
  assign \PCIN[43]  = PCIN[43];
  assign \PCIN[44]  = PCIN[44];
  assign \PCIN[45]  = PCIN[45];
  assign \PCIN[46]  = PCIN[46];
  assign \PCIN[47]  = PCIN[47];
  assign \PCIN[4]  = PCIN[4];
  assign \PCIN[5]  = PCIN[5];
  assign \PCIN[6]  = PCIN[6];
  assign \PCIN[7]  = PCIN[7];
  assign \PCIN[8]  = PCIN[8];
  assign \PCIN[9]  = PCIN[9];
  assign PCOUT[47] = \PCOUT[47] ;
  assign PCOUT[46] = \PCOUT[46] ;
  assign PCOUT[45] = \PCOUT[45] ;
  assign PCOUT[44] = \PCOUT[44] ;
  assign PCOUT[43] = \PCOUT[43] ;
  assign PCOUT[42] = \PCOUT[42] ;
  assign PCOUT[41] = \PCOUT[41] ;
  assign PCOUT[40] = \PCOUT[40] ;
  assign PCOUT[39] = \PCOUT[39] ;
  assign PCOUT[38] = \PCOUT[38] ;
  assign PCOUT[37] = \PCOUT[37] ;
  assign PCOUT[36] = \PCOUT[36] ;
  assign PCOUT[35] = \PCOUT[35] ;
  assign PCOUT[34] = \PCOUT[34] ;
  assign PCOUT[33] = \PCOUT[33] ;
  assign PCOUT[32] = \PCOUT[32] ;
  assign PCOUT[31] = \PCOUT[31] ;
  assign PCOUT[30] = \PCOUT[30] ;
  assign PCOUT[29] = \PCOUT[29] ;
  assign PCOUT[28] = \PCOUT[28] ;
  assign PCOUT[27] = \PCOUT[27] ;
  assign PCOUT[26] = \PCOUT[26] ;
  assign PCOUT[25] = \PCOUT[25] ;
  assign PCOUT[24] = \PCOUT[24] ;
  assign PCOUT[23] = \PCOUT[23] ;
  assign PCOUT[22] = \PCOUT[22] ;
  assign PCOUT[21] = \PCOUT[21] ;
  assign PCOUT[20] = \PCOUT[20] ;
  assign PCOUT[19] = \PCOUT[19] ;
  assign PCOUT[18] = \PCOUT[18] ;
  assign PCOUT[17] = \PCOUT[17] ;
  assign PCOUT[16] = \PCOUT[16] ;
  assign PCOUT[15] = \PCOUT[15] ;
  assign PCOUT[14] = \PCOUT[14] ;
  assign PCOUT[13] = \PCOUT[13] ;
  assign PCOUT[12] = \PCOUT[12] ;
  assign PCOUT[11] = \PCOUT[11] ;
  assign PCOUT[10] = \PCOUT[10] ;
  assign PCOUT[9] = \PCOUT[9] ;
  assign PCOUT[8] = \PCOUT[8] ;
  assign PCOUT[7] = \PCOUT[7] ;
  assign PCOUT[6] = \PCOUT[6] ;
  assign PCOUT[5] = \PCOUT[5] ;
  assign PCOUT[4] = \PCOUT[4] ;
  assign PCOUT[3] = \PCOUT[3] ;
  assign PCOUT[2] = \PCOUT[2] ;
  assign PCOUT[1] = \PCOUT[1] ;
  assign PCOUT[0] = \PCOUT[0] ;
  assign XOROUT[7] = \XOROUT[7] ;
  assign XOROUT[6] = \XOROUT[6] ;
  assign XOROUT[5] = \XOROUT[5] ;
  assign XOROUT[4] = \XOROUT[4] ;
  assign XOROUT[3] = \XOROUT[3] ;
  assign XOROUT[2] = \XOROUT[2] ;
  assign XOROUT[1] = \XOROUT[1] ;
  assign XOROUT[0] = \XOROUT[0] ;
  DSP_ALU #(
    .ALUMODEREG(0),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_OPMODE_INVERTED(9'b000000000),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .MREG(0),
    .OPMODEREG(0),
    .RND(48'h000000000000),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")) 
    DSP_ALU_INST
       (.ALUMODE({\ALUMODE[3] ,\ALUMODE[2] ,\ALUMODE[1] ,\ALUMODE[0] }),
        .ALUMODE10(\DSP_ALU.ALUMODE10 ),
        .ALU_OUT({\DSP_ALU.ALU_OUT<47> ,\DSP_ALU.ALU_OUT<46> ,\DSP_ALU.ALU_OUT<45> ,\DSP_ALU.ALU_OUT<44> ,\DSP_ALU.ALU_OUT<43> ,\DSP_ALU.ALU_OUT<42> ,\DSP_ALU.ALU_OUT<41> ,\DSP_ALU.ALU_OUT<40> ,\DSP_ALU.ALU_OUT<39> ,\DSP_ALU.ALU_OUT<38> ,\DSP_ALU.ALU_OUT<37> ,\DSP_ALU.ALU_OUT<36> ,\DSP_ALU.ALU_OUT<35> ,\DSP_ALU.ALU_OUT<34> ,\DSP_ALU.ALU_OUT<33> ,\DSP_ALU.ALU_OUT<32> ,\DSP_ALU.ALU_OUT<31> ,\DSP_ALU.ALU_OUT<30> ,\DSP_ALU.ALU_OUT<29> ,\DSP_ALU.ALU_OUT<28> ,\DSP_ALU.ALU_OUT<27> ,\DSP_ALU.ALU_OUT<26> ,\DSP_ALU.ALU_OUT<25> ,\DSP_ALU.ALU_OUT<24> ,\DSP_ALU.ALU_OUT<23> ,\DSP_ALU.ALU_OUT<22> ,\DSP_ALU.ALU_OUT<21> ,\DSP_ALU.ALU_OUT<20> ,\DSP_ALU.ALU_OUT<19> ,\DSP_ALU.ALU_OUT<18> ,\DSP_ALU.ALU_OUT<17> ,\DSP_ALU.ALU_OUT<16> ,\DSP_ALU.ALU_OUT<15> ,\DSP_ALU.ALU_OUT<14> ,\DSP_ALU.ALU_OUT<13> ,\DSP_ALU.ALU_OUT<12> ,\DSP_ALU.ALU_OUT<11> ,\DSP_ALU.ALU_OUT<10> ,\DSP_ALU.ALU_OUT<9> ,\DSP_ALU.ALU_OUT<8> ,\DSP_ALU.ALU_OUT<7> ,\DSP_ALU.ALU_OUT<6> ,\DSP_ALU.ALU_OUT<5> ,\DSP_ALU.ALU_OUT<4> ,\DSP_ALU.ALU_OUT<3> ,\DSP_ALU.ALU_OUT<2> ,\DSP_ALU.ALU_OUT<1> ,\DSP_ALU.ALU_OUT<0> }),
        .AMULT26(\DSP_MULTIPLIER.AMULT26 ),
        .A_ALU({\DSP_A_B_DATA.A_ALU<29> ,\DSP_A_B_DATA.A_ALU<28> ,\DSP_A_B_DATA.A_ALU<27> ,\DSP_A_B_DATA.A_ALU<26> ,\DSP_A_B_DATA.A_ALU<25> ,\DSP_A_B_DATA.A_ALU<24> ,\DSP_A_B_DATA.A_ALU<23> ,\DSP_A_B_DATA.A_ALU<22> ,\DSP_A_B_DATA.A_ALU<21> ,\DSP_A_B_DATA.A_ALU<20> ,\DSP_A_B_DATA.A_ALU<19> ,\DSP_A_B_DATA.A_ALU<18> ,\DSP_A_B_DATA.A_ALU<17> ,\DSP_A_B_DATA.A_ALU<16> ,\DSP_A_B_DATA.A_ALU<15> ,\DSP_A_B_DATA.A_ALU<14> ,\DSP_A_B_DATA.A_ALU<13> ,\DSP_A_B_DATA.A_ALU<12> ,\DSP_A_B_DATA.A_ALU<11> ,\DSP_A_B_DATA.A_ALU<10> ,\DSP_A_B_DATA.A_ALU<9> ,\DSP_A_B_DATA.A_ALU<8> ,\DSP_A_B_DATA.A_ALU<7> ,\DSP_A_B_DATA.A_ALU<6> ,\DSP_A_B_DATA.A_ALU<5> ,\DSP_A_B_DATA.A_ALU<4> ,\DSP_A_B_DATA.A_ALU<3> ,\DSP_A_B_DATA.A_ALU<2> ,\DSP_A_B_DATA.A_ALU<1> ,\DSP_A_B_DATA.A_ALU<0> }),
        .BMULT17(\DSP_MULTIPLIER.BMULT17 ),
        .B_ALU({\DSP_A_B_DATA.B_ALU<17> ,\DSP_A_B_DATA.B_ALU<16> ,\DSP_A_B_DATA.B_ALU<15> ,\DSP_A_B_DATA.B_ALU<14> ,\DSP_A_B_DATA.B_ALU<13> ,\DSP_A_B_DATA.B_ALU<12> ,\DSP_A_B_DATA.B_ALU<11> ,\DSP_A_B_DATA.B_ALU<10> ,\DSP_A_B_DATA.B_ALU<9> ,\DSP_A_B_DATA.B_ALU<8> ,\DSP_A_B_DATA.B_ALU<7> ,\DSP_A_B_DATA.B_ALU<6> ,\DSP_A_B_DATA.B_ALU<5> ,\DSP_A_B_DATA.B_ALU<4> ,\DSP_A_B_DATA.B_ALU<3> ,\DSP_A_B_DATA.B_ALU<2> ,\DSP_A_B_DATA.B_ALU<1> ,\DSP_A_B_DATA.B_ALU<0> }),
        .CARRYCASCIN(CARRYCASCIN),
        .CARRYIN(CARRYIN),
        .CARRYINSEL({\CARRYINSEL[2] ,\CARRYINSEL[1] ,\CARRYINSEL[0] }),
        .CCOUT(\DSP_OUTPUT.CCOUT_FB ),
        .CEALUMODE(CEALUMODE),
        .CECARRYIN(CECARRYIN),
        .CECTRL(CECTRL),
        .CEM(CEM),
        .CLK(CLK),
        .COUT({\DSP_ALU.COUT<3> ,\DSP_ALU.COUT<2> ,\DSP_ALU.COUT<1> ,\DSP_ALU.COUT<0> }),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .MULTSIGNIN(MULTSIGNIN),
        .MULTSIGN_ALU(\DSP_ALU.MULTSIGN_ALU ),
        .OPMODE({\OPMODE[8] ,\OPMODE[7] ,\OPMODE[6] ,\OPMODE[5] ,\OPMODE[4] ,\OPMODE[3] ,\OPMODE[2] ,\OPMODE[1] ,\OPMODE[0] }),
        .PCIN({\PCIN[47] ,\PCIN[46] ,\PCIN[45] ,\PCIN[44] ,\PCIN[43] ,\PCIN[42] ,\PCIN[41] ,\PCIN[40] ,\PCIN[39] ,\PCIN[38] ,\PCIN[37] ,\PCIN[36] ,\PCIN[35] ,\PCIN[34] ,\PCIN[33] ,\PCIN[32] ,\PCIN[31] ,\PCIN[30] ,\PCIN[29] ,\PCIN[28] ,\PCIN[27] ,\PCIN[26] ,\PCIN[25] ,\PCIN[24] ,\PCIN[23] ,\PCIN[22] ,\PCIN[21] ,\PCIN[20] ,\PCIN[19] ,\PCIN[18] ,\PCIN[17] ,\PCIN[16] ,\PCIN[15] ,\PCIN[14] ,\PCIN[13] ,\PCIN[12] ,\PCIN[11] ,\PCIN[10] ,\PCIN[9] ,\PCIN[8] ,\PCIN[7] ,\PCIN[6] ,\PCIN[5] ,\PCIN[4] ,\PCIN[3] ,\PCIN[2] ,\PCIN[1] ,\PCIN[0] }),
        .P_FDBK({\DSP_OUTPUT.P_FDBK<47> ,\DSP_OUTPUT.P_FDBK<46> ,\DSP_OUTPUT.P_FDBK<45> ,\DSP_OUTPUT.P_FDBK<44> ,\DSP_OUTPUT.P_FDBK<43> ,\DSP_OUTPUT.P_FDBK<42> ,\DSP_OUTPUT.P_FDBK<41> ,\DSP_OUTPUT.P_FDBK<40> ,\DSP_OUTPUT.P_FDBK<39> ,\DSP_OUTPUT.P_FDBK<38> ,\DSP_OUTPUT.P_FDBK<37> ,\DSP_OUTPUT.P_FDBK<36> ,\DSP_OUTPUT.P_FDBK<35> ,\DSP_OUTPUT.P_FDBK<34> ,\DSP_OUTPUT.P_FDBK<33> ,\DSP_OUTPUT.P_FDBK<32> ,\DSP_OUTPUT.P_FDBK<31> ,\DSP_OUTPUT.P_FDBK<30> ,\DSP_OUTPUT.P_FDBK<29> ,\DSP_OUTPUT.P_FDBK<28> ,\DSP_OUTPUT.P_FDBK<27> ,\DSP_OUTPUT.P_FDBK<26> ,\DSP_OUTPUT.P_FDBK<25> ,\DSP_OUTPUT.P_FDBK<24> ,\DSP_OUTPUT.P_FDBK<23> ,\DSP_OUTPUT.P_FDBK<22> ,\DSP_OUTPUT.P_FDBK<21> ,\DSP_OUTPUT.P_FDBK<20> ,\DSP_OUTPUT.P_FDBK<19> ,\DSP_OUTPUT.P_FDBK<18> ,\DSP_OUTPUT.P_FDBK<17> ,\DSP_OUTPUT.P_FDBK<16> ,\DSP_OUTPUT.P_FDBK<15> ,\DSP_OUTPUT.P_FDBK<14> ,\DSP_OUTPUT.P_FDBK<13> ,\DSP_OUTPUT.P_FDBK<12> ,\DSP_OUTPUT.P_FDBK<11> ,\DSP_OUTPUT.P_FDBK<10> ,\DSP_OUTPUT.P_FDBK<9> ,\DSP_OUTPUT.P_FDBK<8> ,\DSP_OUTPUT.P_FDBK<7> ,\DSP_OUTPUT.P_FDBK<6> ,\DSP_OUTPUT.P_FDBK<5> ,\DSP_OUTPUT.P_FDBK<4> ,\DSP_OUTPUT.P_FDBK<3> ,\DSP_OUTPUT.P_FDBK<2> ,\DSP_OUTPUT.P_FDBK<1> ,\DSP_OUTPUT.P_FDBK<0> }),
        .P_FDBK_47(\DSP_OUTPUT.P_FDBK_47 ),
        .RSTALLCARRYIN(RSTALLCARRYIN),
        .RSTALUMODE(RSTALUMODE),
        .RSTCTRL(RSTCTRL),
        .U_DATA({\DSP_M_DATA.U_DATA<44> ,\DSP_M_DATA.U_DATA<43> ,\DSP_M_DATA.U_DATA<42> ,\DSP_M_DATA.U_DATA<41> ,\DSP_M_DATA.U_DATA<40> ,\DSP_M_DATA.U_DATA<39> ,\DSP_M_DATA.U_DATA<38> ,\DSP_M_DATA.U_DATA<37> ,\DSP_M_DATA.U_DATA<36> ,\DSP_M_DATA.U_DATA<35> ,\DSP_M_DATA.U_DATA<34> ,\DSP_M_DATA.U_DATA<33> ,\DSP_M_DATA.U_DATA<32> ,\DSP_M_DATA.U_DATA<31> ,\DSP_M_DATA.U_DATA<30> ,\DSP_M_DATA.U_DATA<29> ,\DSP_M_DATA.U_DATA<28> ,\DSP_M_DATA.U_DATA<27> ,\DSP_M_DATA.U_DATA<26> ,\DSP_M_DATA.U_DATA<25> ,\DSP_M_DATA.U_DATA<24> ,\DSP_M_DATA.U_DATA<23> ,\DSP_M_DATA.U_DATA<22> ,\DSP_M_DATA.U_DATA<21> ,\DSP_M_DATA.U_DATA<20> ,\DSP_M_DATA.U_DATA<19> ,\DSP_M_DATA.U_DATA<18> ,\DSP_M_DATA.U_DATA<17> ,\DSP_M_DATA.U_DATA<16> ,\DSP_M_DATA.U_DATA<15> ,\DSP_M_DATA.U_DATA<14> ,\DSP_M_DATA.U_DATA<13> ,\DSP_M_DATA.U_DATA<12> ,\DSP_M_DATA.U_DATA<11> ,\DSP_M_DATA.U_DATA<10> ,\DSP_M_DATA.U_DATA<9> ,\DSP_M_DATA.U_DATA<8> ,\DSP_M_DATA.U_DATA<7> ,\DSP_M_DATA.U_DATA<6> ,\DSP_M_DATA.U_DATA<5> ,\DSP_M_DATA.U_DATA<4> ,\DSP_M_DATA.U_DATA<3> ,\DSP_M_DATA.U_DATA<2> ,\DSP_M_DATA.U_DATA<1> ,\DSP_M_DATA.U_DATA<0> }),
        .V_DATA({\DSP_M_DATA.V_DATA<44> ,\DSP_M_DATA.V_DATA<43> ,\DSP_M_DATA.V_DATA<42> ,\DSP_M_DATA.V_DATA<41> ,\DSP_M_DATA.V_DATA<40> ,\DSP_M_DATA.V_DATA<39> ,\DSP_M_DATA.V_DATA<38> ,\DSP_M_DATA.V_DATA<37> ,\DSP_M_DATA.V_DATA<36> ,\DSP_M_DATA.V_DATA<35> ,\DSP_M_DATA.V_DATA<34> ,\DSP_M_DATA.V_DATA<33> ,\DSP_M_DATA.V_DATA<32> ,\DSP_M_DATA.V_DATA<31> ,\DSP_M_DATA.V_DATA<30> ,\DSP_M_DATA.V_DATA<29> ,\DSP_M_DATA.V_DATA<28> ,\DSP_M_DATA.V_DATA<27> ,\DSP_M_DATA.V_DATA<26> ,\DSP_M_DATA.V_DATA<25> ,\DSP_M_DATA.V_DATA<24> ,\DSP_M_DATA.V_DATA<23> ,\DSP_M_DATA.V_DATA<22> ,\DSP_M_DATA.V_DATA<21> ,\DSP_M_DATA.V_DATA<20> ,\DSP_M_DATA.V_DATA<19> ,\DSP_M_DATA.V_DATA<18> ,\DSP_M_DATA.V_DATA<17> ,\DSP_M_DATA.V_DATA<16> ,\DSP_M_DATA.V_DATA<15> ,\DSP_M_DATA.V_DATA<14> ,\DSP_M_DATA.V_DATA<13> ,\DSP_M_DATA.V_DATA<12> ,\DSP_M_DATA.V_DATA<11> ,\DSP_M_DATA.V_DATA<10> ,\DSP_M_DATA.V_DATA<9> ,\DSP_M_DATA.V_DATA<8> ,\DSP_M_DATA.V_DATA<7> ,\DSP_M_DATA.V_DATA<6> ,\DSP_M_DATA.V_DATA<5> ,\DSP_M_DATA.V_DATA<4> ,\DSP_M_DATA.V_DATA<3> ,\DSP_M_DATA.V_DATA<2> ,\DSP_M_DATA.V_DATA<1> ,\DSP_M_DATA.V_DATA<0> }),
        .XOR_MX({\DSP_ALU.XOR_MX<7> ,\DSP_ALU.XOR_MX<6> ,\DSP_ALU.XOR_MX<5> ,\DSP_ALU.XOR_MX<4> ,\DSP_ALU.XOR_MX<3> ,\DSP_ALU.XOR_MX<2> ,\DSP_ALU.XOR_MX<1> ,\DSP_ALU.XOR_MX<0> }));
  DSP_A_B_DATA #(
    .ACASCREG(0),
    .AREG(0),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0)) 
    DSP_A_B_DATA_INST
       (.A({\A[29] ,\A[28] ,\A[27] ,\A[26] ,\A[25] ,\A[24] ,\A[23] ,\A[22] ,\A[21] ,\A[20] ,\A[19] ,\A[18] ,\A[17] ,\A[16] ,\A[15] ,\A[14] ,\A[13] ,\A[12] ,\A[11] ,\A[10] ,\A[9] ,\A[8] ,\A[7] ,\A[6] ,\A[5] ,\A[4] ,\A[3] ,\A[2] ,\A[1] ,\A[0] }),
        .A1_DATA({\DSP_A_B_DATA.A1_DATA<26> ,\DSP_A_B_DATA.A1_DATA<25> ,\DSP_A_B_DATA.A1_DATA<24> ,\DSP_A_B_DATA.A1_DATA<23> ,\DSP_A_B_DATA.A1_DATA<22> ,\DSP_A_B_DATA.A1_DATA<21> ,\DSP_A_B_DATA.A1_DATA<20> ,\DSP_A_B_DATA.A1_DATA<19> ,\DSP_A_B_DATA.A1_DATA<18> ,\DSP_A_B_DATA.A1_DATA<17> ,\DSP_A_B_DATA.A1_DATA<16> ,\DSP_A_B_DATA.A1_DATA<15> ,\DSP_A_B_DATA.A1_DATA<14> ,\DSP_A_B_DATA.A1_DATA<13> ,\DSP_A_B_DATA.A1_DATA<12> ,\DSP_A_B_DATA.A1_DATA<11> ,\DSP_A_B_DATA.A1_DATA<10> ,\DSP_A_B_DATA.A1_DATA<9> ,\DSP_A_B_DATA.A1_DATA<8> ,\DSP_A_B_DATA.A1_DATA<7> ,\DSP_A_B_DATA.A1_DATA<6> ,\DSP_A_B_DATA.A1_DATA<5> ,\DSP_A_B_DATA.A1_DATA<4> ,\DSP_A_B_DATA.A1_DATA<3> ,\DSP_A_B_DATA.A1_DATA<2> ,\DSP_A_B_DATA.A1_DATA<1> ,\DSP_A_B_DATA.A1_DATA<0> }),
        .A2_DATA({\DSP_A_B_DATA.A2_DATA<26> ,\DSP_A_B_DATA.A2_DATA<25> ,\DSP_A_B_DATA.A2_DATA<24> ,\DSP_A_B_DATA.A2_DATA<23> ,\DSP_A_B_DATA.A2_DATA<22> ,\DSP_A_B_DATA.A2_DATA<21> ,\DSP_A_B_DATA.A2_DATA<20> ,\DSP_A_B_DATA.A2_DATA<19> ,\DSP_A_B_DATA.A2_DATA<18> ,\DSP_A_B_DATA.A2_DATA<17> ,\DSP_A_B_DATA.A2_DATA<16> ,\DSP_A_B_DATA.A2_DATA<15> ,\DSP_A_B_DATA.A2_DATA<14> ,\DSP_A_B_DATA.A2_DATA<13> ,\DSP_A_B_DATA.A2_DATA<12> ,\DSP_A_B_DATA.A2_DATA<11> ,\DSP_A_B_DATA.A2_DATA<10> ,\DSP_A_B_DATA.A2_DATA<9> ,\DSP_A_B_DATA.A2_DATA<8> ,\DSP_A_B_DATA.A2_DATA<7> ,\DSP_A_B_DATA.A2_DATA<6> ,\DSP_A_B_DATA.A2_DATA<5> ,\DSP_A_B_DATA.A2_DATA<4> ,\DSP_A_B_DATA.A2_DATA<3> ,\DSP_A_B_DATA.A2_DATA<2> ,\DSP_A_B_DATA.A2_DATA<1> ,\DSP_A_B_DATA.A2_DATA<0> }),
        .ACIN({\ACIN[29] ,\ACIN[28] ,\ACIN[27] ,\ACIN[26] ,\ACIN[25] ,\ACIN[24] ,\ACIN[23] ,\ACIN[22] ,\ACIN[21] ,\ACIN[20] ,\ACIN[19] ,\ACIN[18] ,\ACIN[17] ,\ACIN[16] ,\ACIN[15] ,\ACIN[14] ,\ACIN[13] ,\ACIN[12] ,\ACIN[11] ,\ACIN[10] ,\ACIN[9] ,\ACIN[8] ,\ACIN[7] ,\ACIN[6] ,\ACIN[5] ,\ACIN[4] ,\ACIN[3] ,\ACIN[2] ,\ACIN[1] ,\ACIN[0] }),
        .ACOUT({\ACOUT[29] ,\ACOUT[28] ,\ACOUT[27] ,\ACOUT[26] ,\ACOUT[25] ,\ACOUT[24] ,\ACOUT[23] ,\ACOUT[22] ,\ACOUT[21] ,\ACOUT[20] ,\ACOUT[19] ,\ACOUT[18] ,\ACOUT[17] ,\ACOUT[16] ,\ACOUT[15] ,\ACOUT[14] ,\ACOUT[13] ,\ACOUT[12] ,\ACOUT[11] ,\ACOUT[10] ,\ACOUT[9] ,\ACOUT[8] ,\ACOUT[7] ,\ACOUT[6] ,\ACOUT[5] ,\ACOUT[4] ,\ACOUT[3] ,\ACOUT[2] ,\ACOUT[1] ,\ACOUT[0] }),
        .A_ALU({\DSP_A_B_DATA.A_ALU<29> ,\DSP_A_B_DATA.A_ALU<28> ,\DSP_A_B_DATA.A_ALU<27> ,\DSP_A_B_DATA.A_ALU<26> ,\DSP_A_B_DATA.A_ALU<25> ,\DSP_A_B_DATA.A_ALU<24> ,\DSP_A_B_DATA.A_ALU<23> ,\DSP_A_B_DATA.A_ALU<22> ,\DSP_A_B_DATA.A_ALU<21> ,\DSP_A_B_DATA.A_ALU<20> ,\DSP_A_B_DATA.A_ALU<19> ,\DSP_A_B_DATA.A_ALU<18> ,\DSP_A_B_DATA.A_ALU<17> ,\DSP_A_B_DATA.A_ALU<16> ,\DSP_A_B_DATA.A_ALU<15> ,\DSP_A_B_DATA.A_ALU<14> ,\DSP_A_B_DATA.A_ALU<13> ,\DSP_A_B_DATA.A_ALU<12> ,\DSP_A_B_DATA.A_ALU<11> ,\DSP_A_B_DATA.A_ALU<10> ,\DSP_A_B_DATA.A_ALU<9> ,\DSP_A_B_DATA.A_ALU<8> ,\DSP_A_B_DATA.A_ALU<7> ,\DSP_A_B_DATA.A_ALU<6> ,\DSP_A_B_DATA.A_ALU<5> ,\DSP_A_B_DATA.A_ALU<4> ,\DSP_A_B_DATA.A_ALU<3> ,\DSP_A_B_DATA.A_ALU<2> ,\DSP_A_B_DATA.A_ALU<1> ,\DSP_A_B_DATA.A_ALU<0> }),
        .B({\B[17] ,\B[16] ,\B[15] ,\B[14] ,\B[13] ,\B[12] ,\B[11] ,\B[10] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,\B[0] }),
        .B1_DATA({\DSP_A_B_DATA.B1_DATA<17> ,\DSP_A_B_DATA.B1_DATA<16> ,\DSP_A_B_DATA.B1_DATA<15> ,\DSP_A_B_DATA.B1_DATA<14> ,\DSP_A_B_DATA.B1_DATA<13> ,\DSP_A_B_DATA.B1_DATA<12> ,\DSP_A_B_DATA.B1_DATA<11> ,\DSP_A_B_DATA.B1_DATA<10> ,\DSP_A_B_DATA.B1_DATA<9> ,\DSP_A_B_DATA.B1_DATA<8> ,\DSP_A_B_DATA.B1_DATA<7> ,\DSP_A_B_DATA.B1_DATA<6> ,\DSP_A_B_DATA.B1_DATA<5> ,\DSP_A_B_DATA.B1_DATA<4> ,\DSP_A_B_DATA.B1_DATA<3> ,\DSP_A_B_DATA.B1_DATA<2> ,\DSP_A_B_DATA.B1_DATA<1> ,\DSP_A_B_DATA.B1_DATA<0> }),
        .B2_DATA({\DSP_A_B_DATA.B2_DATA<17> ,\DSP_A_B_DATA.B2_DATA<16> ,\DSP_A_B_DATA.B2_DATA<15> ,\DSP_A_B_DATA.B2_DATA<14> ,\DSP_A_B_DATA.B2_DATA<13> ,\DSP_A_B_DATA.B2_DATA<12> ,\DSP_A_B_DATA.B2_DATA<11> ,\DSP_A_B_DATA.B2_DATA<10> ,\DSP_A_B_DATA.B2_DATA<9> ,\DSP_A_B_DATA.B2_DATA<8> ,\DSP_A_B_DATA.B2_DATA<7> ,\DSP_A_B_DATA.B2_DATA<6> ,\DSP_A_B_DATA.B2_DATA<5> ,\DSP_A_B_DATA.B2_DATA<4> ,\DSP_A_B_DATA.B2_DATA<3> ,\DSP_A_B_DATA.B2_DATA<2> ,\DSP_A_B_DATA.B2_DATA<1> ,\DSP_A_B_DATA.B2_DATA<0> }),
        .BCIN({\BCIN[17] ,\BCIN[16] ,\BCIN[15] ,\BCIN[14] ,\BCIN[13] ,\BCIN[12] ,\BCIN[11] ,\BCIN[10] ,\BCIN[9] ,\BCIN[8] ,\BCIN[7] ,\BCIN[6] ,\BCIN[5] ,\BCIN[4] ,\BCIN[3] ,\BCIN[2] ,\BCIN[1] ,\BCIN[0] }),
        .BCOUT({\BCOUT[17] ,\BCOUT[16] ,\BCOUT[15] ,\BCOUT[14] ,\BCOUT[13] ,\BCOUT[12] ,\BCOUT[11] ,\BCOUT[10] ,\BCOUT[9] ,\BCOUT[8] ,\BCOUT[7] ,\BCOUT[6] ,\BCOUT[5] ,\BCOUT[4] ,\BCOUT[3] ,\BCOUT[2] ,\BCOUT[1] ,\BCOUT[0] }),
        .B_ALU({\DSP_A_B_DATA.B_ALU<17> ,\DSP_A_B_DATA.B_ALU<16> ,\DSP_A_B_DATA.B_ALU<15> ,\DSP_A_B_DATA.B_ALU<14> ,\DSP_A_B_DATA.B_ALU<13> ,\DSP_A_B_DATA.B_ALU<12> ,\DSP_A_B_DATA.B_ALU<11> ,\DSP_A_B_DATA.B_ALU<10> ,\DSP_A_B_DATA.B_ALU<9> ,\DSP_A_B_DATA.B_ALU<8> ,\DSP_A_B_DATA.B_ALU<7> ,\DSP_A_B_DATA.B_ALU<6> ,\DSP_A_B_DATA.B_ALU<5> ,\DSP_A_B_DATA.B_ALU<4> ,\DSP_A_B_DATA.B_ALU<3> ,\DSP_A_B_DATA.B_ALU<2> ,\DSP_A_B_DATA.B_ALU<1> ,\DSP_A_B_DATA.B_ALU<0> }),
        .CEA1(CEA1),
        .CEA2(CEA2),
        .CEB1(CEB1),
        .CEB2(CEB2),
        .CLK(CLK),
        .RSTA(RSTA),
        .RSTB(RSTB));
  DSP_C_DATA #(
    .CREG(0),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0)) 
    DSP_C_DATA_INST
       (.C({\C[47] ,\C[46] ,\C[45] ,\C[44] ,\C[43] ,\C[42] ,\C[41] ,\C[40] ,\C[39] ,\C[38] ,\C[37] ,\C[36] ,\C[35] ,\C[34] ,\C[33] ,\C[32] ,\C[31] ,\C[30] ,\C[29] ,\C[28] ,\C[27] ,\C[26] ,\C[25] ,\C[24] ,\C[23] ,\C[22] ,\C[21] ,\C[20] ,\C[19] ,\C[18] ,\C[17] ,\C[16] ,\C[15] ,\C[14] ,\C[13] ,\C[12] ,\C[11] ,\C[10] ,\C[9] ,\C[8] ,\C[7] ,\C[6] ,\C[5] ,\C[4] ,\C[3] ,\C[2] ,\C[1] ,\C[0] }),
        .CEC(CEC),
        .CLK(CLK),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .RSTC(RSTC));
  DSP_MULTIPLIER #(
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .USE_MULT("MULTIPLY")) 
    DSP_MULTIPLIER_INST
       (.A2A1({\DSP_PREADD_DATA.A2A1<26> ,\DSP_PREADD_DATA.A2A1<25> ,\DSP_PREADD_DATA.A2A1<24> ,\DSP_PREADD_DATA.A2A1<23> ,\DSP_PREADD_DATA.A2A1<22> ,\DSP_PREADD_DATA.A2A1<21> ,\DSP_PREADD_DATA.A2A1<20> ,\DSP_PREADD_DATA.A2A1<19> ,\DSP_PREADD_DATA.A2A1<18> ,\DSP_PREADD_DATA.A2A1<17> ,\DSP_PREADD_DATA.A2A1<16> ,\DSP_PREADD_DATA.A2A1<15> ,\DSP_PREADD_DATA.A2A1<14> ,\DSP_PREADD_DATA.A2A1<13> ,\DSP_PREADD_DATA.A2A1<12> ,\DSP_PREADD_DATA.A2A1<11> ,\DSP_PREADD_DATA.A2A1<10> ,\DSP_PREADD_DATA.A2A1<9> ,\DSP_PREADD_DATA.A2A1<8> ,\DSP_PREADD_DATA.A2A1<7> ,\DSP_PREADD_DATA.A2A1<6> ,\DSP_PREADD_DATA.A2A1<5> ,\DSP_PREADD_DATA.A2A1<4> ,\DSP_PREADD_DATA.A2A1<3> ,\DSP_PREADD_DATA.A2A1<2> ,\DSP_PREADD_DATA.A2A1<1> ,\DSP_PREADD_DATA.A2A1<0> }),
        .AD_DATA({\DSP_PREADD_DATA.AD_DATA<26> ,\DSP_PREADD_DATA.AD_DATA<25> ,\DSP_PREADD_DATA.AD_DATA<24> ,\DSP_PREADD_DATA.AD_DATA<23> ,\DSP_PREADD_DATA.AD_DATA<22> ,\DSP_PREADD_DATA.AD_DATA<21> ,\DSP_PREADD_DATA.AD_DATA<20> ,\DSP_PREADD_DATA.AD_DATA<19> ,\DSP_PREADD_DATA.AD_DATA<18> ,\DSP_PREADD_DATA.AD_DATA<17> ,\DSP_PREADD_DATA.AD_DATA<16> ,\DSP_PREADD_DATA.AD_DATA<15> ,\DSP_PREADD_DATA.AD_DATA<14> ,\DSP_PREADD_DATA.AD_DATA<13> ,\DSP_PREADD_DATA.AD_DATA<12> ,\DSP_PREADD_DATA.AD_DATA<11> ,\DSP_PREADD_DATA.AD_DATA<10> ,\DSP_PREADD_DATA.AD_DATA<9> ,\DSP_PREADD_DATA.AD_DATA<8> ,\DSP_PREADD_DATA.AD_DATA<7> ,\DSP_PREADD_DATA.AD_DATA<6> ,\DSP_PREADD_DATA.AD_DATA<5> ,\DSP_PREADD_DATA.AD_DATA<4> ,\DSP_PREADD_DATA.AD_DATA<3> ,\DSP_PREADD_DATA.AD_DATA<2> ,\DSP_PREADD_DATA.AD_DATA<1> ,\DSP_PREADD_DATA.AD_DATA<0> }),
        .AMULT26(\DSP_MULTIPLIER.AMULT26 ),
        .B2B1({\DSP_PREADD_DATA.B2B1<17> ,\DSP_PREADD_DATA.B2B1<16> ,\DSP_PREADD_DATA.B2B1<15> ,\DSP_PREADD_DATA.B2B1<14> ,\DSP_PREADD_DATA.B2B1<13> ,\DSP_PREADD_DATA.B2B1<12> ,\DSP_PREADD_DATA.B2B1<11> ,\DSP_PREADD_DATA.B2B1<10> ,\DSP_PREADD_DATA.B2B1<9> ,\DSP_PREADD_DATA.B2B1<8> ,\DSP_PREADD_DATA.B2B1<7> ,\DSP_PREADD_DATA.B2B1<6> ,\DSP_PREADD_DATA.B2B1<5> ,\DSP_PREADD_DATA.B2B1<4> ,\DSP_PREADD_DATA.B2B1<3> ,\DSP_PREADD_DATA.B2B1<2> ,\DSP_PREADD_DATA.B2B1<1> ,\DSP_PREADD_DATA.B2B1<0> }),
        .BMULT17(\DSP_MULTIPLIER.BMULT17 ),
        .U({\DSP_MULTIPLIER.U<44> ,\DSP_MULTIPLIER.U<43> ,\DSP_MULTIPLIER.U<42> ,\DSP_MULTIPLIER.U<41> ,\DSP_MULTIPLIER.U<40> ,\DSP_MULTIPLIER.U<39> ,\DSP_MULTIPLIER.U<38> ,\DSP_MULTIPLIER.U<37> ,\DSP_MULTIPLIER.U<36> ,\DSP_MULTIPLIER.U<35> ,\DSP_MULTIPLIER.U<34> ,\DSP_MULTIPLIER.U<33> ,\DSP_MULTIPLIER.U<32> ,\DSP_MULTIPLIER.U<31> ,\DSP_MULTIPLIER.U<30> ,\DSP_MULTIPLIER.U<29> ,\DSP_MULTIPLIER.U<28> ,\DSP_MULTIPLIER.U<27> ,\DSP_MULTIPLIER.U<26> ,\DSP_MULTIPLIER.U<25> ,\DSP_MULTIPLIER.U<24> ,\DSP_MULTIPLIER.U<23> ,\DSP_MULTIPLIER.U<22> ,\DSP_MULTIPLIER.U<21> ,\DSP_MULTIPLIER.U<20> ,\DSP_MULTIPLIER.U<19> ,\DSP_MULTIPLIER.U<18> ,\DSP_MULTIPLIER.U<17> ,\DSP_MULTIPLIER.U<16> ,\DSP_MULTIPLIER.U<15> ,\DSP_MULTIPLIER.U<14> ,\DSP_MULTIPLIER.U<13> ,\DSP_MULTIPLIER.U<12> ,\DSP_MULTIPLIER.U<11> ,\DSP_MULTIPLIER.U<10> ,\DSP_MULTIPLIER.U<9> ,\DSP_MULTIPLIER.U<8> ,\DSP_MULTIPLIER.U<7> ,\DSP_MULTIPLIER.U<6> ,\DSP_MULTIPLIER.U<5> ,\DSP_MULTIPLIER.U<4> ,\DSP_MULTIPLIER.U<3> ,\DSP_MULTIPLIER.U<2> ,\DSP_MULTIPLIER.U<1> ,\DSP_MULTIPLIER.U<0> }),
        .V({\DSP_MULTIPLIER.V<44> ,\DSP_MULTIPLIER.V<43> ,\DSP_MULTIPLIER.V<42> ,\DSP_MULTIPLIER.V<41> ,\DSP_MULTIPLIER.V<40> ,\DSP_MULTIPLIER.V<39> ,\DSP_MULTIPLIER.V<38> ,\DSP_MULTIPLIER.V<37> ,\DSP_MULTIPLIER.V<36> ,\DSP_MULTIPLIER.V<35> ,\DSP_MULTIPLIER.V<34> ,\DSP_MULTIPLIER.V<33> ,\DSP_MULTIPLIER.V<32> ,\DSP_MULTIPLIER.V<31> ,\DSP_MULTIPLIER.V<30> ,\DSP_MULTIPLIER.V<29> ,\DSP_MULTIPLIER.V<28> ,\DSP_MULTIPLIER.V<27> ,\DSP_MULTIPLIER.V<26> ,\DSP_MULTIPLIER.V<25> ,\DSP_MULTIPLIER.V<24> ,\DSP_MULTIPLIER.V<23> ,\DSP_MULTIPLIER.V<22> ,\DSP_MULTIPLIER.V<21> ,\DSP_MULTIPLIER.V<20> ,\DSP_MULTIPLIER.V<19> ,\DSP_MULTIPLIER.V<18> ,\DSP_MULTIPLIER.V<17> ,\DSP_MULTIPLIER.V<16> ,\DSP_MULTIPLIER.V<15> ,\DSP_MULTIPLIER.V<14> ,\DSP_MULTIPLIER.V<13> ,\DSP_MULTIPLIER.V<12> ,\DSP_MULTIPLIER.V<11> ,\DSP_MULTIPLIER.V<10> ,\DSP_MULTIPLIER.V<9> ,\DSP_MULTIPLIER.V<8> ,\DSP_MULTIPLIER.V<7> ,\DSP_MULTIPLIER.V<6> ,\DSP_MULTIPLIER.V<5> ,\DSP_MULTIPLIER.V<4> ,\DSP_MULTIPLIER.V<3> ,\DSP_MULTIPLIER.V<2> ,\DSP_MULTIPLIER.V<1> ,\DSP_MULTIPLIER.V<0> }));
  DSP_M_DATA #(
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .MREG(0)) 
    DSP_M_DATA_INST
       (.CEM(CEM),
        .CLK(CLK),
        .RSTM(RSTM),
        .U({\DSP_MULTIPLIER.U<44> ,\DSP_MULTIPLIER.U<43> ,\DSP_MULTIPLIER.U<42> ,\DSP_MULTIPLIER.U<41> ,\DSP_MULTIPLIER.U<40> ,\DSP_MULTIPLIER.U<39> ,\DSP_MULTIPLIER.U<38> ,\DSP_MULTIPLIER.U<37> ,\DSP_MULTIPLIER.U<36> ,\DSP_MULTIPLIER.U<35> ,\DSP_MULTIPLIER.U<34> ,\DSP_MULTIPLIER.U<33> ,\DSP_MULTIPLIER.U<32> ,\DSP_MULTIPLIER.U<31> ,\DSP_MULTIPLIER.U<30> ,\DSP_MULTIPLIER.U<29> ,\DSP_MULTIPLIER.U<28> ,\DSP_MULTIPLIER.U<27> ,\DSP_MULTIPLIER.U<26> ,\DSP_MULTIPLIER.U<25> ,\DSP_MULTIPLIER.U<24> ,\DSP_MULTIPLIER.U<23> ,\DSP_MULTIPLIER.U<22> ,\DSP_MULTIPLIER.U<21> ,\DSP_MULTIPLIER.U<20> ,\DSP_MULTIPLIER.U<19> ,\DSP_MULTIPLIER.U<18> ,\DSP_MULTIPLIER.U<17> ,\DSP_MULTIPLIER.U<16> ,\DSP_MULTIPLIER.U<15> ,\DSP_MULTIPLIER.U<14> ,\DSP_MULTIPLIER.U<13> ,\DSP_MULTIPLIER.U<12> ,\DSP_MULTIPLIER.U<11> ,\DSP_MULTIPLIER.U<10> ,\DSP_MULTIPLIER.U<9> ,\DSP_MULTIPLIER.U<8> ,\DSP_MULTIPLIER.U<7> ,\DSP_MULTIPLIER.U<6> ,\DSP_MULTIPLIER.U<5> ,\DSP_MULTIPLIER.U<4> ,\DSP_MULTIPLIER.U<3> ,\DSP_MULTIPLIER.U<2> ,\DSP_MULTIPLIER.U<1> ,\DSP_MULTIPLIER.U<0> }),
        .U_DATA({\DSP_M_DATA.U_DATA<44> ,\DSP_M_DATA.U_DATA<43> ,\DSP_M_DATA.U_DATA<42> ,\DSP_M_DATA.U_DATA<41> ,\DSP_M_DATA.U_DATA<40> ,\DSP_M_DATA.U_DATA<39> ,\DSP_M_DATA.U_DATA<38> ,\DSP_M_DATA.U_DATA<37> ,\DSP_M_DATA.U_DATA<36> ,\DSP_M_DATA.U_DATA<35> ,\DSP_M_DATA.U_DATA<34> ,\DSP_M_DATA.U_DATA<33> ,\DSP_M_DATA.U_DATA<32> ,\DSP_M_DATA.U_DATA<31> ,\DSP_M_DATA.U_DATA<30> ,\DSP_M_DATA.U_DATA<29> ,\DSP_M_DATA.U_DATA<28> ,\DSP_M_DATA.U_DATA<27> ,\DSP_M_DATA.U_DATA<26> ,\DSP_M_DATA.U_DATA<25> ,\DSP_M_DATA.U_DATA<24> ,\DSP_M_DATA.U_DATA<23> ,\DSP_M_DATA.U_DATA<22> ,\DSP_M_DATA.U_DATA<21> ,\DSP_M_DATA.U_DATA<20> ,\DSP_M_DATA.U_DATA<19> ,\DSP_M_DATA.U_DATA<18> ,\DSP_M_DATA.U_DATA<17> ,\DSP_M_DATA.U_DATA<16> ,\DSP_M_DATA.U_DATA<15> ,\DSP_M_DATA.U_DATA<14> ,\DSP_M_DATA.U_DATA<13> ,\DSP_M_DATA.U_DATA<12> ,\DSP_M_DATA.U_DATA<11> ,\DSP_M_DATA.U_DATA<10> ,\DSP_M_DATA.U_DATA<9> ,\DSP_M_DATA.U_DATA<8> ,\DSP_M_DATA.U_DATA<7> ,\DSP_M_DATA.U_DATA<6> ,\DSP_M_DATA.U_DATA<5> ,\DSP_M_DATA.U_DATA<4> ,\DSP_M_DATA.U_DATA<3> ,\DSP_M_DATA.U_DATA<2> ,\DSP_M_DATA.U_DATA<1> ,\DSP_M_DATA.U_DATA<0> }),
        .V({\DSP_MULTIPLIER.V<44> ,\DSP_MULTIPLIER.V<43> ,\DSP_MULTIPLIER.V<42> ,\DSP_MULTIPLIER.V<41> ,\DSP_MULTIPLIER.V<40> ,\DSP_MULTIPLIER.V<39> ,\DSP_MULTIPLIER.V<38> ,\DSP_MULTIPLIER.V<37> ,\DSP_MULTIPLIER.V<36> ,\DSP_MULTIPLIER.V<35> ,\DSP_MULTIPLIER.V<34> ,\DSP_MULTIPLIER.V<33> ,\DSP_MULTIPLIER.V<32> ,\DSP_MULTIPLIER.V<31> ,\DSP_MULTIPLIER.V<30> ,\DSP_MULTIPLIER.V<29> ,\DSP_MULTIPLIER.V<28> ,\DSP_MULTIPLIER.V<27> ,\DSP_MULTIPLIER.V<26> ,\DSP_MULTIPLIER.V<25> ,\DSP_MULTIPLIER.V<24> ,\DSP_MULTIPLIER.V<23> ,\DSP_MULTIPLIER.V<22> ,\DSP_MULTIPLIER.V<21> ,\DSP_MULTIPLIER.V<20> ,\DSP_MULTIPLIER.V<19> ,\DSP_MULTIPLIER.V<18> ,\DSP_MULTIPLIER.V<17> ,\DSP_MULTIPLIER.V<16> ,\DSP_MULTIPLIER.V<15> ,\DSP_MULTIPLIER.V<14> ,\DSP_MULTIPLIER.V<13> ,\DSP_MULTIPLIER.V<12> ,\DSP_MULTIPLIER.V<11> ,\DSP_MULTIPLIER.V<10> ,\DSP_MULTIPLIER.V<9> ,\DSP_MULTIPLIER.V<8> ,\DSP_MULTIPLIER.V<7> ,\DSP_MULTIPLIER.V<6> ,\DSP_MULTIPLIER.V<5> ,\DSP_MULTIPLIER.V<4> ,\DSP_MULTIPLIER.V<3> ,\DSP_MULTIPLIER.V<2> ,\DSP_MULTIPLIER.V<1> ,\DSP_MULTIPLIER.V<0> }),
        .V_DATA({\DSP_M_DATA.V_DATA<44> ,\DSP_M_DATA.V_DATA<43> ,\DSP_M_DATA.V_DATA<42> ,\DSP_M_DATA.V_DATA<41> ,\DSP_M_DATA.V_DATA<40> ,\DSP_M_DATA.V_DATA<39> ,\DSP_M_DATA.V_DATA<38> ,\DSP_M_DATA.V_DATA<37> ,\DSP_M_DATA.V_DATA<36> ,\DSP_M_DATA.V_DATA<35> ,\DSP_M_DATA.V_DATA<34> ,\DSP_M_DATA.V_DATA<33> ,\DSP_M_DATA.V_DATA<32> ,\DSP_M_DATA.V_DATA<31> ,\DSP_M_DATA.V_DATA<30> ,\DSP_M_DATA.V_DATA<29> ,\DSP_M_DATA.V_DATA<28> ,\DSP_M_DATA.V_DATA<27> ,\DSP_M_DATA.V_DATA<26> ,\DSP_M_DATA.V_DATA<25> ,\DSP_M_DATA.V_DATA<24> ,\DSP_M_DATA.V_DATA<23> ,\DSP_M_DATA.V_DATA<22> ,\DSP_M_DATA.V_DATA<21> ,\DSP_M_DATA.V_DATA<20> ,\DSP_M_DATA.V_DATA<19> ,\DSP_M_DATA.V_DATA<18> ,\DSP_M_DATA.V_DATA<17> ,\DSP_M_DATA.V_DATA<16> ,\DSP_M_DATA.V_DATA<15> ,\DSP_M_DATA.V_DATA<14> ,\DSP_M_DATA.V_DATA<13> ,\DSP_M_DATA.V_DATA<12> ,\DSP_M_DATA.V_DATA<11> ,\DSP_M_DATA.V_DATA<10> ,\DSP_M_DATA.V_DATA<9> ,\DSP_M_DATA.V_DATA<8> ,\DSP_M_DATA.V_DATA<7> ,\DSP_M_DATA.V_DATA<6> ,\DSP_M_DATA.V_DATA<5> ,\DSP_M_DATA.V_DATA<4> ,\DSP_M_DATA.V_DATA<3> ,\DSP_M_DATA.V_DATA<2> ,\DSP_M_DATA.V_DATA<1> ,\DSP_M_DATA.V_DATA<0> }));
  DSP_OUTPUT #(
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h3FFFFFFFFFFF),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_PATTERN_DETECT("NO_PATDET")) 
    DSP_OUTPUT_INST
       (.ALUMODE10(\DSP_ALU.ALUMODE10 ),
        .ALU_OUT({\DSP_ALU.ALU_OUT<47> ,\DSP_ALU.ALU_OUT<46> ,\DSP_ALU.ALU_OUT<45> ,\DSP_ALU.ALU_OUT<44> ,\DSP_ALU.ALU_OUT<43> ,\DSP_ALU.ALU_OUT<42> ,\DSP_ALU.ALU_OUT<41> ,\DSP_ALU.ALU_OUT<40> ,\DSP_ALU.ALU_OUT<39> ,\DSP_ALU.ALU_OUT<38> ,\DSP_ALU.ALU_OUT<37> ,\DSP_ALU.ALU_OUT<36> ,\DSP_ALU.ALU_OUT<35> ,\DSP_ALU.ALU_OUT<34> ,\DSP_ALU.ALU_OUT<33> ,\DSP_ALU.ALU_OUT<32> ,\DSP_ALU.ALU_OUT<31> ,\DSP_ALU.ALU_OUT<30> ,\DSP_ALU.ALU_OUT<29> ,\DSP_ALU.ALU_OUT<28> ,\DSP_ALU.ALU_OUT<27> ,\DSP_ALU.ALU_OUT<26> ,\DSP_ALU.ALU_OUT<25> ,\DSP_ALU.ALU_OUT<24> ,\DSP_ALU.ALU_OUT<23> ,\DSP_ALU.ALU_OUT<22> ,\DSP_ALU.ALU_OUT<21> ,\DSP_ALU.ALU_OUT<20> ,\DSP_ALU.ALU_OUT<19> ,\DSP_ALU.ALU_OUT<18> ,\DSP_ALU.ALU_OUT<17> ,\DSP_ALU.ALU_OUT<16> ,\DSP_ALU.ALU_OUT<15> ,\DSP_ALU.ALU_OUT<14> ,\DSP_ALU.ALU_OUT<13> ,\DSP_ALU.ALU_OUT<12> ,\DSP_ALU.ALU_OUT<11> ,\DSP_ALU.ALU_OUT<10> ,\DSP_ALU.ALU_OUT<9> ,\DSP_ALU.ALU_OUT<8> ,\DSP_ALU.ALU_OUT<7> ,\DSP_ALU.ALU_OUT<6> ,\DSP_ALU.ALU_OUT<5> ,\DSP_ALU.ALU_OUT<4> ,\DSP_ALU.ALU_OUT<3> ,\DSP_ALU.ALU_OUT<2> ,\DSP_ALU.ALU_OUT<1> ,\DSP_ALU.ALU_OUT<0> }),
        .CARRYCASCOUT(CARRYCASCOUT),
        .CARRYOUT({\CARRYOUT[3] ,\CARRYOUT[2] ,\CARRYOUT[1] ,\CARRYOUT[0] }),
        .CCOUT_FB(\DSP_OUTPUT.CCOUT_FB ),
        .CEP(CEP),
        .CLK(CLK),
        .COUT({\DSP_ALU.COUT<3> ,\DSP_ALU.COUT<2> ,\DSP_ALU.COUT<1> ,\DSP_ALU.COUT<0> }),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .MULTSIGNOUT(MULTSIGNOUT),
        .MULTSIGN_ALU(\DSP_ALU.MULTSIGN_ALU ),
        .OVERFLOW(OVERFLOW),
        .P({\P[47] ,\P[46] ,\P[45] ,\P[44] ,\P[43] ,\P[42] ,\P[41] ,\P[40] ,\P[39] ,\P[38] ,\P[37] ,\P[36] ,\P[35] ,\P[34] ,\P[33] ,\P[32] ,\P[31] ,\P[30] ,\P[29] ,\P[28] ,\P[27] ,\P[26] ,\P[25] ,\P[24] ,\P[23] ,\P[22] ,\P[21] ,\P[20] ,\P[19] ,\P[18] ,\P[17] ,\P[16] ,\P[15] ,\P[14] ,\P[13] ,\P[12] ,\P[11] ,\P[10] ,\P[9] ,\P[8] ,\P[7] ,\P[6] ,\P[5] ,\P[4] ,\P[3] ,\P[2] ,\P[1] ,\P[0] }),
        .PATTERN_B_DETECT(PATTERNBDETECT),
        .PATTERN_DETECT(PATTERNDETECT),
        .PCOUT({\PCOUT[47] ,\PCOUT[46] ,\PCOUT[45] ,\PCOUT[44] ,\PCOUT[43] ,\PCOUT[42] ,\PCOUT[41] ,\PCOUT[40] ,\PCOUT[39] ,\PCOUT[38] ,\PCOUT[37] ,\PCOUT[36] ,\PCOUT[35] ,\PCOUT[34] ,\PCOUT[33] ,\PCOUT[32] ,\PCOUT[31] ,\PCOUT[30] ,\PCOUT[29] ,\PCOUT[28] ,\PCOUT[27] ,\PCOUT[26] ,\PCOUT[25] ,\PCOUT[24] ,\PCOUT[23] ,\PCOUT[22] ,\PCOUT[21] ,\PCOUT[20] ,\PCOUT[19] ,\PCOUT[18] ,\PCOUT[17] ,\PCOUT[16] ,\PCOUT[15] ,\PCOUT[14] ,\PCOUT[13] ,\PCOUT[12] ,\PCOUT[11] ,\PCOUT[10] ,\PCOUT[9] ,\PCOUT[8] ,\PCOUT[7] ,\PCOUT[6] ,\PCOUT[5] ,\PCOUT[4] ,\PCOUT[3] ,\PCOUT[2] ,\PCOUT[1] ,\PCOUT[0] }),
        .P_FDBK({\DSP_OUTPUT.P_FDBK<47> ,\DSP_OUTPUT.P_FDBK<46> ,\DSP_OUTPUT.P_FDBK<45> ,\DSP_OUTPUT.P_FDBK<44> ,\DSP_OUTPUT.P_FDBK<43> ,\DSP_OUTPUT.P_FDBK<42> ,\DSP_OUTPUT.P_FDBK<41> ,\DSP_OUTPUT.P_FDBK<40> ,\DSP_OUTPUT.P_FDBK<39> ,\DSP_OUTPUT.P_FDBK<38> ,\DSP_OUTPUT.P_FDBK<37> ,\DSP_OUTPUT.P_FDBK<36> ,\DSP_OUTPUT.P_FDBK<35> ,\DSP_OUTPUT.P_FDBK<34> ,\DSP_OUTPUT.P_FDBK<33> ,\DSP_OUTPUT.P_FDBK<32> ,\DSP_OUTPUT.P_FDBK<31> ,\DSP_OUTPUT.P_FDBK<30> ,\DSP_OUTPUT.P_FDBK<29> ,\DSP_OUTPUT.P_FDBK<28> ,\DSP_OUTPUT.P_FDBK<27> ,\DSP_OUTPUT.P_FDBK<26> ,\DSP_OUTPUT.P_FDBK<25> ,\DSP_OUTPUT.P_FDBK<24> ,\DSP_OUTPUT.P_FDBK<23> ,\DSP_OUTPUT.P_FDBK<22> ,\DSP_OUTPUT.P_FDBK<21> ,\DSP_OUTPUT.P_FDBK<20> ,\DSP_OUTPUT.P_FDBK<19> ,\DSP_OUTPUT.P_FDBK<18> ,\DSP_OUTPUT.P_FDBK<17> ,\DSP_OUTPUT.P_FDBK<16> ,\DSP_OUTPUT.P_FDBK<15> ,\DSP_OUTPUT.P_FDBK<14> ,\DSP_OUTPUT.P_FDBK<13> ,\DSP_OUTPUT.P_FDBK<12> ,\DSP_OUTPUT.P_FDBK<11> ,\DSP_OUTPUT.P_FDBK<10> ,\DSP_OUTPUT.P_FDBK<9> ,\DSP_OUTPUT.P_FDBK<8> ,\DSP_OUTPUT.P_FDBK<7> ,\DSP_OUTPUT.P_FDBK<6> ,\DSP_OUTPUT.P_FDBK<5> ,\DSP_OUTPUT.P_FDBK<4> ,\DSP_OUTPUT.P_FDBK<3> ,\DSP_OUTPUT.P_FDBK<2> ,\DSP_OUTPUT.P_FDBK<1> ,\DSP_OUTPUT.P_FDBK<0> }),
        .P_FDBK_47(\DSP_OUTPUT.P_FDBK_47 ),
        .RSTP(RSTP),
        .UNDERFLOW(UNDERFLOW),
        .XOROUT({\XOROUT[7] ,\XOROUT[6] ,\XOROUT[5] ,\XOROUT[4] ,\XOROUT[3] ,\XOROUT[2] ,\XOROUT[1] ,\XOROUT[0] }),
        .XOR_MX({\DSP_ALU.XOR_MX<7> ,\DSP_ALU.XOR_MX<6> ,\DSP_ALU.XOR_MX<5> ,\DSP_ALU.XOR_MX<4> ,\DSP_ALU.XOR_MX<3> ,\DSP_ALU.XOR_MX<2> ,\DSP_ALU.XOR_MX<1> ,\DSP_ALU.XOR_MX<0> }));
  DSP_PREADD_DATA #(
    .ADREG(1),
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .DREG(1),
    .INMODEREG(0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .PREADDINSEL("A"),
    .USE_MULT("MULTIPLY")) 
    DSP_PREADD_DATA_INST
       (.A1_DATA({\DSP_A_B_DATA.A1_DATA<26> ,\DSP_A_B_DATA.A1_DATA<25> ,\DSP_A_B_DATA.A1_DATA<24> ,\DSP_A_B_DATA.A1_DATA<23> ,\DSP_A_B_DATA.A1_DATA<22> ,\DSP_A_B_DATA.A1_DATA<21> ,\DSP_A_B_DATA.A1_DATA<20> ,\DSP_A_B_DATA.A1_DATA<19> ,\DSP_A_B_DATA.A1_DATA<18> ,\DSP_A_B_DATA.A1_DATA<17> ,\DSP_A_B_DATA.A1_DATA<16> ,\DSP_A_B_DATA.A1_DATA<15> ,\DSP_A_B_DATA.A1_DATA<14> ,\DSP_A_B_DATA.A1_DATA<13> ,\DSP_A_B_DATA.A1_DATA<12> ,\DSP_A_B_DATA.A1_DATA<11> ,\DSP_A_B_DATA.A1_DATA<10> ,\DSP_A_B_DATA.A1_DATA<9> ,\DSP_A_B_DATA.A1_DATA<8> ,\DSP_A_B_DATA.A1_DATA<7> ,\DSP_A_B_DATA.A1_DATA<6> ,\DSP_A_B_DATA.A1_DATA<5> ,\DSP_A_B_DATA.A1_DATA<4> ,\DSP_A_B_DATA.A1_DATA<3> ,\DSP_A_B_DATA.A1_DATA<2> ,\DSP_A_B_DATA.A1_DATA<1> ,\DSP_A_B_DATA.A1_DATA<0> }),
        .A2A1({\DSP_PREADD_DATA.A2A1<26> ,\DSP_PREADD_DATA.A2A1<25> ,\DSP_PREADD_DATA.A2A1<24> ,\DSP_PREADD_DATA.A2A1<23> ,\DSP_PREADD_DATA.A2A1<22> ,\DSP_PREADD_DATA.A2A1<21> ,\DSP_PREADD_DATA.A2A1<20> ,\DSP_PREADD_DATA.A2A1<19> ,\DSP_PREADD_DATA.A2A1<18> ,\DSP_PREADD_DATA.A2A1<17> ,\DSP_PREADD_DATA.A2A1<16> ,\DSP_PREADD_DATA.A2A1<15> ,\DSP_PREADD_DATA.A2A1<14> ,\DSP_PREADD_DATA.A2A1<13> ,\DSP_PREADD_DATA.A2A1<12> ,\DSP_PREADD_DATA.A2A1<11> ,\DSP_PREADD_DATA.A2A1<10> ,\DSP_PREADD_DATA.A2A1<9> ,\DSP_PREADD_DATA.A2A1<8> ,\DSP_PREADD_DATA.A2A1<7> ,\DSP_PREADD_DATA.A2A1<6> ,\DSP_PREADD_DATA.A2A1<5> ,\DSP_PREADD_DATA.A2A1<4> ,\DSP_PREADD_DATA.A2A1<3> ,\DSP_PREADD_DATA.A2A1<2> ,\DSP_PREADD_DATA.A2A1<1> ,\DSP_PREADD_DATA.A2A1<0> }),
        .A2_DATA({\DSP_A_B_DATA.A2_DATA<26> ,\DSP_A_B_DATA.A2_DATA<25> ,\DSP_A_B_DATA.A2_DATA<24> ,\DSP_A_B_DATA.A2_DATA<23> ,\DSP_A_B_DATA.A2_DATA<22> ,\DSP_A_B_DATA.A2_DATA<21> ,\DSP_A_B_DATA.A2_DATA<20> ,\DSP_A_B_DATA.A2_DATA<19> ,\DSP_A_B_DATA.A2_DATA<18> ,\DSP_A_B_DATA.A2_DATA<17> ,\DSP_A_B_DATA.A2_DATA<16> ,\DSP_A_B_DATA.A2_DATA<15> ,\DSP_A_B_DATA.A2_DATA<14> ,\DSP_A_B_DATA.A2_DATA<13> ,\DSP_A_B_DATA.A2_DATA<12> ,\DSP_A_B_DATA.A2_DATA<11> ,\DSP_A_B_DATA.A2_DATA<10> ,\DSP_A_B_DATA.A2_DATA<9> ,\DSP_A_B_DATA.A2_DATA<8> ,\DSP_A_B_DATA.A2_DATA<7> ,\DSP_A_B_DATA.A2_DATA<6> ,\DSP_A_B_DATA.A2_DATA<5> ,\DSP_A_B_DATA.A2_DATA<4> ,\DSP_A_B_DATA.A2_DATA<3> ,\DSP_A_B_DATA.A2_DATA<2> ,\DSP_A_B_DATA.A2_DATA<1> ,\DSP_A_B_DATA.A2_DATA<0> }),
        .AD({\DSP_PREADD.AD<26> ,\DSP_PREADD.AD<25> ,\DSP_PREADD.AD<24> ,\DSP_PREADD.AD<23> ,\DSP_PREADD.AD<22> ,\DSP_PREADD.AD<21> ,\DSP_PREADD.AD<20> ,\DSP_PREADD.AD<19> ,\DSP_PREADD.AD<18> ,\DSP_PREADD.AD<17> ,\DSP_PREADD.AD<16> ,\DSP_PREADD.AD<15> ,\DSP_PREADD.AD<14> ,\DSP_PREADD.AD<13> ,\DSP_PREADD.AD<12> ,\DSP_PREADD.AD<11> ,\DSP_PREADD.AD<10> ,\DSP_PREADD.AD<9> ,\DSP_PREADD.AD<8> ,\DSP_PREADD.AD<7> ,\DSP_PREADD.AD<6> ,\DSP_PREADD.AD<5> ,\DSP_PREADD.AD<4> ,\DSP_PREADD.AD<3> ,\DSP_PREADD.AD<2> ,\DSP_PREADD.AD<1> ,\DSP_PREADD.AD<0> }),
        .ADDSUB(\DSP_PREADD_DATA.ADDSUB ),
        .AD_DATA({\DSP_PREADD_DATA.AD_DATA<26> ,\DSP_PREADD_DATA.AD_DATA<25> ,\DSP_PREADD_DATA.AD_DATA<24> ,\DSP_PREADD_DATA.AD_DATA<23> ,\DSP_PREADD_DATA.AD_DATA<22> ,\DSP_PREADD_DATA.AD_DATA<21> ,\DSP_PREADD_DATA.AD_DATA<20> ,\DSP_PREADD_DATA.AD_DATA<19> ,\DSP_PREADD_DATA.AD_DATA<18> ,\DSP_PREADD_DATA.AD_DATA<17> ,\DSP_PREADD_DATA.AD_DATA<16> ,\DSP_PREADD_DATA.AD_DATA<15> ,\DSP_PREADD_DATA.AD_DATA<14> ,\DSP_PREADD_DATA.AD_DATA<13> ,\DSP_PREADD_DATA.AD_DATA<12> ,\DSP_PREADD_DATA.AD_DATA<11> ,\DSP_PREADD_DATA.AD_DATA<10> ,\DSP_PREADD_DATA.AD_DATA<9> ,\DSP_PREADD_DATA.AD_DATA<8> ,\DSP_PREADD_DATA.AD_DATA<7> ,\DSP_PREADD_DATA.AD_DATA<6> ,\DSP_PREADD_DATA.AD_DATA<5> ,\DSP_PREADD_DATA.AD_DATA<4> ,\DSP_PREADD_DATA.AD_DATA<3> ,\DSP_PREADD_DATA.AD_DATA<2> ,\DSP_PREADD_DATA.AD_DATA<1> ,\DSP_PREADD_DATA.AD_DATA<0> }),
        .B1_DATA({\DSP_A_B_DATA.B1_DATA<17> ,\DSP_A_B_DATA.B1_DATA<16> ,\DSP_A_B_DATA.B1_DATA<15> ,\DSP_A_B_DATA.B1_DATA<14> ,\DSP_A_B_DATA.B1_DATA<13> ,\DSP_A_B_DATA.B1_DATA<12> ,\DSP_A_B_DATA.B1_DATA<11> ,\DSP_A_B_DATA.B1_DATA<10> ,\DSP_A_B_DATA.B1_DATA<9> ,\DSP_A_B_DATA.B1_DATA<8> ,\DSP_A_B_DATA.B1_DATA<7> ,\DSP_A_B_DATA.B1_DATA<6> ,\DSP_A_B_DATA.B1_DATA<5> ,\DSP_A_B_DATA.B1_DATA<4> ,\DSP_A_B_DATA.B1_DATA<3> ,\DSP_A_B_DATA.B1_DATA<2> ,\DSP_A_B_DATA.B1_DATA<1> ,\DSP_A_B_DATA.B1_DATA<0> }),
        .B2B1({\DSP_PREADD_DATA.B2B1<17> ,\DSP_PREADD_DATA.B2B1<16> ,\DSP_PREADD_DATA.B2B1<15> ,\DSP_PREADD_DATA.B2B1<14> ,\DSP_PREADD_DATA.B2B1<13> ,\DSP_PREADD_DATA.B2B1<12> ,\DSP_PREADD_DATA.B2B1<11> ,\DSP_PREADD_DATA.B2B1<10> ,\DSP_PREADD_DATA.B2B1<9> ,\DSP_PREADD_DATA.B2B1<8> ,\DSP_PREADD_DATA.B2B1<7> ,\DSP_PREADD_DATA.B2B1<6> ,\DSP_PREADD_DATA.B2B1<5> ,\DSP_PREADD_DATA.B2B1<4> ,\DSP_PREADD_DATA.B2B1<3> ,\DSP_PREADD_DATA.B2B1<2> ,\DSP_PREADD_DATA.B2B1<1> ,\DSP_PREADD_DATA.B2B1<0> }),
        .B2_DATA({\DSP_A_B_DATA.B2_DATA<17> ,\DSP_A_B_DATA.B2_DATA<16> ,\DSP_A_B_DATA.B2_DATA<15> ,\DSP_A_B_DATA.B2_DATA<14> ,\DSP_A_B_DATA.B2_DATA<13> ,\DSP_A_B_DATA.B2_DATA<12> ,\DSP_A_B_DATA.B2_DATA<11> ,\DSP_A_B_DATA.B2_DATA<10> ,\DSP_A_B_DATA.B2_DATA<9> ,\DSP_A_B_DATA.B2_DATA<8> ,\DSP_A_B_DATA.B2_DATA<7> ,\DSP_A_B_DATA.B2_DATA<6> ,\DSP_A_B_DATA.B2_DATA<5> ,\DSP_A_B_DATA.B2_DATA<4> ,\DSP_A_B_DATA.B2_DATA<3> ,\DSP_A_B_DATA.B2_DATA<2> ,\DSP_A_B_DATA.B2_DATA<1> ,\DSP_A_B_DATA.B2_DATA<0> }),
        .CEAD(CEAD),
        .CED(CED),
        .CEINMODE(CEINMODE),
        .CLK(CLK),
        .DIN({\D[26] ,\D[25] ,\D[24] ,\D[23] ,\D[22] ,\D[21] ,\D[20] ,\D[19] ,\D[18] ,\D[17] ,\D[16] ,\D[15] ,\D[14] ,\D[13] ,\D[12] ,\D[11] ,\D[10] ,\D[9] ,\D[8] ,\D[7] ,\D[6] ,\D[5] ,\D[4] ,\D[3] ,\D[2] ,\D[1] ,\D[0] }),
        .D_DATA({\DSP_PREADD_DATA.D_DATA<26> ,\DSP_PREADD_DATA.D_DATA<25> ,\DSP_PREADD_DATA.D_DATA<24> ,\DSP_PREADD_DATA.D_DATA<23> ,\DSP_PREADD_DATA.D_DATA<22> ,\DSP_PREADD_DATA.D_DATA<21> ,\DSP_PREADD_DATA.D_DATA<20> ,\DSP_PREADD_DATA.D_DATA<19> ,\DSP_PREADD_DATA.D_DATA<18> ,\DSP_PREADD_DATA.D_DATA<17> ,\DSP_PREADD_DATA.D_DATA<16> ,\DSP_PREADD_DATA.D_DATA<15> ,\DSP_PREADD_DATA.D_DATA<14> ,\DSP_PREADD_DATA.D_DATA<13> ,\DSP_PREADD_DATA.D_DATA<12> ,\DSP_PREADD_DATA.D_DATA<11> ,\DSP_PREADD_DATA.D_DATA<10> ,\DSP_PREADD_DATA.D_DATA<9> ,\DSP_PREADD_DATA.D_DATA<8> ,\DSP_PREADD_DATA.D_DATA<7> ,\DSP_PREADD_DATA.D_DATA<6> ,\DSP_PREADD_DATA.D_DATA<5> ,\DSP_PREADD_DATA.D_DATA<4> ,\DSP_PREADD_DATA.D_DATA<3> ,\DSP_PREADD_DATA.D_DATA<2> ,\DSP_PREADD_DATA.D_DATA<1> ,\DSP_PREADD_DATA.D_DATA<0> }),
        .INMODE({\INMODE[4] ,\INMODE[3] ,\INMODE[2] ,\INMODE[1] ,\INMODE[0] }),
        .INMODE_2(\DSP_PREADD_DATA.INMODE_2 ),
        .PREADD_AB({\DSP_PREADD_DATA.PREADD_AB<26> ,\DSP_PREADD_DATA.PREADD_AB<25> ,\DSP_PREADD_DATA.PREADD_AB<24> ,\DSP_PREADD_DATA.PREADD_AB<23> ,\DSP_PREADD_DATA.PREADD_AB<22> ,\DSP_PREADD_DATA.PREADD_AB<21> ,\DSP_PREADD_DATA.PREADD_AB<20> ,\DSP_PREADD_DATA.PREADD_AB<19> ,\DSP_PREADD_DATA.PREADD_AB<18> ,\DSP_PREADD_DATA.PREADD_AB<17> ,\DSP_PREADD_DATA.PREADD_AB<16> ,\DSP_PREADD_DATA.PREADD_AB<15> ,\DSP_PREADD_DATA.PREADD_AB<14> ,\DSP_PREADD_DATA.PREADD_AB<13> ,\DSP_PREADD_DATA.PREADD_AB<12> ,\DSP_PREADD_DATA.PREADD_AB<11> ,\DSP_PREADD_DATA.PREADD_AB<10> ,\DSP_PREADD_DATA.PREADD_AB<9> ,\DSP_PREADD_DATA.PREADD_AB<8> ,\DSP_PREADD_DATA.PREADD_AB<7> ,\DSP_PREADD_DATA.PREADD_AB<6> ,\DSP_PREADD_DATA.PREADD_AB<5> ,\DSP_PREADD_DATA.PREADD_AB<4> ,\DSP_PREADD_DATA.PREADD_AB<3> ,\DSP_PREADD_DATA.PREADD_AB<2> ,\DSP_PREADD_DATA.PREADD_AB<1> ,\DSP_PREADD_DATA.PREADD_AB<0> }),
        .RSTD(RSTD),
        .RSTINMODE(RSTINMODE));
  DSP_PREADD DSP_PREADD_INST
       (.AD({\DSP_PREADD.AD<26> ,\DSP_PREADD.AD<25> ,\DSP_PREADD.AD<24> ,\DSP_PREADD.AD<23> ,\DSP_PREADD.AD<22> ,\DSP_PREADD.AD<21> ,\DSP_PREADD.AD<20> ,\DSP_PREADD.AD<19> ,\DSP_PREADD.AD<18> ,\DSP_PREADD.AD<17> ,\DSP_PREADD.AD<16> ,\DSP_PREADD.AD<15> ,\DSP_PREADD.AD<14> ,\DSP_PREADD.AD<13> ,\DSP_PREADD.AD<12> ,\DSP_PREADD.AD<11> ,\DSP_PREADD.AD<10> ,\DSP_PREADD.AD<9> ,\DSP_PREADD.AD<8> ,\DSP_PREADD.AD<7> ,\DSP_PREADD.AD<6> ,\DSP_PREADD.AD<5> ,\DSP_PREADD.AD<4> ,\DSP_PREADD.AD<3> ,\DSP_PREADD.AD<2> ,\DSP_PREADD.AD<1> ,\DSP_PREADD.AD<0> }),
        .ADDSUB(\DSP_PREADD_DATA.ADDSUB ),
        .D_DATA({\DSP_PREADD_DATA.D_DATA<26> ,\DSP_PREADD_DATA.D_DATA<25> ,\DSP_PREADD_DATA.D_DATA<24> ,\DSP_PREADD_DATA.D_DATA<23> ,\DSP_PREADD_DATA.D_DATA<22> ,\DSP_PREADD_DATA.D_DATA<21> ,\DSP_PREADD_DATA.D_DATA<20> ,\DSP_PREADD_DATA.D_DATA<19> ,\DSP_PREADD_DATA.D_DATA<18> ,\DSP_PREADD_DATA.D_DATA<17> ,\DSP_PREADD_DATA.D_DATA<16> ,\DSP_PREADD_DATA.D_DATA<15> ,\DSP_PREADD_DATA.D_DATA<14> ,\DSP_PREADD_DATA.D_DATA<13> ,\DSP_PREADD_DATA.D_DATA<12> ,\DSP_PREADD_DATA.D_DATA<11> ,\DSP_PREADD_DATA.D_DATA<10> ,\DSP_PREADD_DATA.D_DATA<9> ,\DSP_PREADD_DATA.D_DATA<8> ,\DSP_PREADD_DATA.D_DATA<7> ,\DSP_PREADD_DATA.D_DATA<6> ,\DSP_PREADD_DATA.D_DATA<5> ,\DSP_PREADD_DATA.D_DATA<4> ,\DSP_PREADD_DATA.D_DATA<3> ,\DSP_PREADD_DATA.D_DATA<2> ,\DSP_PREADD_DATA.D_DATA<1> ,\DSP_PREADD_DATA.D_DATA<0> }),
        .INMODE2(\DSP_PREADD_DATA.INMODE_2 ),
        .PREADD_AB({\DSP_PREADD_DATA.PREADD_AB<26> ,\DSP_PREADD_DATA.PREADD_AB<25> ,\DSP_PREADD_DATA.PREADD_AB<24> ,\DSP_PREADD_DATA.PREADD_AB<23> ,\DSP_PREADD_DATA.PREADD_AB<22> ,\DSP_PREADD_DATA.PREADD_AB<21> ,\DSP_PREADD_DATA.PREADD_AB<20> ,\DSP_PREADD_DATA.PREADD_AB<19> ,\DSP_PREADD_DATA.PREADD_AB<18> ,\DSP_PREADD_DATA.PREADD_AB<17> ,\DSP_PREADD_DATA.PREADD_AB<16> ,\DSP_PREADD_DATA.PREADD_AB<15> ,\DSP_PREADD_DATA.PREADD_AB<14> ,\DSP_PREADD_DATA.PREADD_AB<13> ,\DSP_PREADD_DATA.PREADD_AB<12> ,\DSP_PREADD_DATA.PREADD_AB<11> ,\DSP_PREADD_DATA.PREADD_AB<10> ,\DSP_PREADD_DATA.PREADD_AB<9> ,\DSP_PREADD_DATA.PREADD_AB<8> ,\DSP_PREADD_DATA.PREADD_AB<7> ,\DSP_PREADD_DATA.PREADD_AB<6> ,\DSP_PREADD_DATA.PREADD_AB<5> ,\DSP_PREADD_DATA.PREADD_AB<4> ,\DSP_PREADD_DATA.PREADD_AB<3> ,\DSP_PREADD_DATA.PREADD_AB<2> ,\DSP_PREADD_DATA.PREADD_AB<1> ,\DSP_PREADD_DATA.PREADD_AB<0> }));
endmodule

module DSP48E2_HD32741
   (ACOUT,
    BCOUT,
    CARRYCASCOUT,
    CARRYOUT,
    MULTSIGNOUT,
    OVERFLOW,
    PATTERNBDETECT,
    PATTERNDETECT,
    PCOUT,
    P,
    UNDERFLOW,
    XOROUT,
    ACIN,
    ALUMODE,
    A,
    BCIN,
    B,
    CARRYCASCIN,
    CARRYIN,
    CARRYINSEL,
    CEA1,
    CEA2,
    CEAD,
    CEALUMODE,
    CEB1,
    CEB2,
    CEC,
    CECARRYIN,
    CECTRL,
    CED,
    CEINMODE,
    CEM,
    CEP,
    CLK,
    C,
    D,
    INMODE,
    MULTSIGNIN,
    OPMODE,
    PCIN,
    RSTA,
    RSTALLCARRYIN,
    RSTALUMODE,
    RSTB,
    RSTC,
    RSTCTRL,
    RSTD,
    RSTINMODE,
    RSTM,
    RSTP);
  output [29:0]ACOUT;
  output [17:0]BCOUT;
  output CARRYCASCOUT;
  output [3:0]CARRYOUT;
  output MULTSIGNOUT;
  output OVERFLOW;
  output PATTERNBDETECT;
  output PATTERNDETECT;
  output [47:0]PCOUT;
  output [47:0]P;
  output UNDERFLOW;
  output [7:0]XOROUT;
  input [29:0]ACIN;
  input [3:0]ALUMODE;
  input [29:0]A;
  input [17:0]BCIN;
  input [17:0]B;
  input CARRYCASCIN;
  input CARRYIN;
  input [2:0]CARRYINSEL;
  input CEA1;
  input CEA2;
  input CEAD;
  input CEALUMODE;
  input CEB1;
  input CEB2;
  input CEC;
  input CECARRYIN;
  input CECTRL;
  input CED;
  input CEINMODE;
  input CEM;
  input CEP;
  input CLK;
  input [47:0]C;
  input [26:0]D;
  input [4:0]INMODE;
  input MULTSIGNIN;
  input [8:0]OPMODE;
  input [47:0]PCIN;
  input RSTA;
  input RSTALLCARRYIN;
  input RSTALUMODE;
  input RSTB;
  input RSTC;
  input RSTCTRL;
  input RSTD;
  input RSTINMODE;
  input RSTM;
  input RSTP;

  wire \ACIN[0] ;
  wire \ACIN[10] ;
  wire \ACIN[11] ;
  wire \ACIN[12] ;
  wire \ACIN[13] ;
  wire \ACIN[14] ;
  wire \ACIN[15] ;
  wire \ACIN[16] ;
  wire \ACIN[17] ;
  wire \ACIN[18] ;
  wire \ACIN[19] ;
  wire \ACIN[1] ;
  wire \ACIN[20] ;
  wire \ACIN[21] ;
  wire \ACIN[22] ;
  wire \ACIN[23] ;
  wire \ACIN[24] ;
  wire \ACIN[25] ;
  wire \ACIN[26] ;
  wire \ACIN[27] ;
  wire \ACIN[28] ;
  wire \ACIN[29] ;
  wire \ACIN[2] ;
  wire \ACIN[3] ;
  wire \ACIN[4] ;
  wire \ACIN[5] ;
  wire \ACIN[6] ;
  wire \ACIN[7] ;
  wire \ACIN[8] ;
  wire \ACIN[9] ;
  wire \ACOUT[0] ;
  wire \ACOUT[10] ;
  wire \ACOUT[11] ;
  wire \ACOUT[12] ;
  wire \ACOUT[13] ;
  wire \ACOUT[14] ;
  wire \ACOUT[15] ;
  wire \ACOUT[16] ;
  wire \ACOUT[17] ;
  wire \ACOUT[18] ;
  wire \ACOUT[19] ;
  wire \ACOUT[1] ;
  wire \ACOUT[20] ;
  wire \ACOUT[21] ;
  wire \ACOUT[22] ;
  wire \ACOUT[23] ;
  wire \ACOUT[24] ;
  wire \ACOUT[25] ;
  wire \ACOUT[26] ;
  wire \ACOUT[27] ;
  wire \ACOUT[28] ;
  wire \ACOUT[29] ;
  wire \ACOUT[2] ;
  wire \ACOUT[3] ;
  wire \ACOUT[4] ;
  wire \ACOUT[5] ;
  wire \ACOUT[6] ;
  wire \ACOUT[7] ;
  wire \ACOUT[8] ;
  wire \ACOUT[9] ;
  wire \ALUMODE[0] ;
  wire \ALUMODE[1] ;
  wire \ALUMODE[2] ;
  wire \ALUMODE[3] ;
  wire \A[0] ;
  wire \A[10] ;
  wire \A[11] ;
  wire \A[12] ;
  wire \A[13] ;
  wire \A[14] ;
  wire \A[15] ;
  wire \A[16] ;
  wire \A[17] ;
  wire \A[18] ;
  wire \A[19] ;
  wire \A[1] ;
  wire \A[20] ;
  wire \A[21] ;
  wire \A[22] ;
  wire \A[23] ;
  wire \A[24] ;
  wire \A[25] ;
  wire \A[26] ;
  wire \A[27] ;
  wire \A[28] ;
  wire \A[29] ;
  wire \A[2] ;
  wire \A[3] ;
  wire \A[4] ;
  wire \A[5] ;
  wire \A[6] ;
  wire \A[7] ;
  wire \A[8] ;
  wire \A[9] ;
  wire \BCIN[0] ;
  wire \BCIN[10] ;
  wire \BCIN[11] ;
  wire \BCIN[12] ;
  wire \BCIN[13] ;
  wire \BCIN[14] ;
  wire \BCIN[15] ;
  wire \BCIN[16] ;
  wire \BCIN[17] ;
  wire \BCIN[1] ;
  wire \BCIN[2] ;
  wire \BCIN[3] ;
  wire \BCIN[4] ;
  wire \BCIN[5] ;
  wire \BCIN[6] ;
  wire \BCIN[7] ;
  wire \BCIN[8] ;
  wire \BCIN[9] ;
  wire \BCOUT[0] ;
  wire \BCOUT[10] ;
  wire \BCOUT[11] ;
  wire \BCOUT[12] ;
  wire \BCOUT[13] ;
  wire \BCOUT[14] ;
  wire \BCOUT[15] ;
  wire \BCOUT[16] ;
  wire \BCOUT[17] ;
  wire \BCOUT[1] ;
  wire \BCOUT[2] ;
  wire \BCOUT[3] ;
  wire \BCOUT[4] ;
  wire \BCOUT[5] ;
  wire \BCOUT[6] ;
  wire \BCOUT[7] ;
  wire \BCOUT[8] ;
  wire \BCOUT[9] ;
  wire \B[0] ;
  wire \B[10] ;
  wire \B[11] ;
  wire \B[12] ;
  wire \B[13] ;
  wire \B[14] ;
  wire \B[15] ;
  wire \B[16] ;
  wire \B[17] ;
  wire \B[1] ;
  wire \B[2] ;
  wire \B[3] ;
  wire \B[4] ;
  wire \B[5] ;
  wire \B[6] ;
  wire \B[7] ;
  wire \B[8] ;
  wire \B[9] ;
  wire CARRYCASCIN;
  wire CARRYCASCOUT;
  wire CARRYIN;
  wire \CARRYINSEL[0] ;
  wire \CARRYINSEL[1] ;
  wire \CARRYINSEL[2] ;
  wire \CARRYOUT[0] ;
  wire \CARRYOUT[1] ;
  wire \CARRYOUT[2] ;
  wire \CARRYOUT[3] ;
  wire CEA1;
  wire CEA2;
  wire CEAD;
  wire CEALUMODE;
  wire CEB1;
  wire CEB2;
  wire CEC;
  wire CECARRYIN;
  wire CECTRL;
  wire CED;
  wire CEINMODE;
  wire CEM;
  wire CEP;
  wire CLK;
  wire \C[0] ;
  wire \C[10] ;
  wire \C[11] ;
  wire \C[12] ;
  wire \C[13] ;
  wire \C[14] ;
  wire \C[15] ;
  wire \C[16] ;
  wire \C[17] ;
  wire \C[18] ;
  wire \C[19] ;
  wire \C[1] ;
  wire \C[20] ;
  wire \C[21] ;
  wire \C[22] ;
  wire \C[23] ;
  wire \C[24] ;
  wire \C[25] ;
  wire \C[26] ;
  wire \C[27] ;
  wire \C[28] ;
  wire \C[29] ;
  wire \C[2] ;
  wire \C[30] ;
  wire \C[31] ;
  wire \C[32] ;
  wire \C[33] ;
  wire \C[34] ;
  wire \C[35] ;
  wire \C[36] ;
  wire \C[37] ;
  wire \C[38] ;
  wire \C[39] ;
  wire \C[3] ;
  wire \C[40] ;
  wire \C[41] ;
  wire \C[42] ;
  wire \C[43] ;
  wire \C[44] ;
  wire \C[45] ;
  wire \C[46] ;
  wire \C[47] ;
  wire \C[4] ;
  wire \C[5] ;
  wire \C[6] ;
  wire \C[7] ;
  wire \C[8] ;
  wire \C[9] ;
  wire \DSP_ALU.ALUMODE10 ;
  wire \DSP_ALU.ALU_OUT<0> ;
  wire \DSP_ALU.ALU_OUT<10> ;
  wire \DSP_ALU.ALU_OUT<11> ;
  wire \DSP_ALU.ALU_OUT<12> ;
  wire \DSP_ALU.ALU_OUT<13> ;
  wire \DSP_ALU.ALU_OUT<14> ;
  wire \DSP_ALU.ALU_OUT<15> ;
  wire \DSP_ALU.ALU_OUT<16> ;
  wire \DSP_ALU.ALU_OUT<17> ;
  wire \DSP_ALU.ALU_OUT<18> ;
  wire \DSP_ALU.ALU_OUT<19> ;
  wire \DSP_ALU.ALU_OUT<1> ;
  wire \DSP_ALU.ALU_OUT<20> ;
  wire \DSP_ALU.ALU_OUT<21> ;
  wire \DSP_ALU.ALU_OUT<22> ;
  wire \DSP_ALU.ALU_OUT<23> ;
  wire \DSP_ALU.ALU_OUT<24> ;
  wire \DSP_ALU.ALU_OUT<25> ;
  wire \DSP_ALU.ALU_OUT<26> ;
  wire \DSP_ALU.ALU_OUT<27> ;
  wire \DSP_ALU.ALU_OUT<28> ;
  wire \DSP_ALU.ALU_OUT<29> ;
  wire \DSP_ALU.ALU_OUT<2> ;
  wire \DSP_ALU.ALU_OUT<30> ;
  wire \DSP_ALU.ALU_OUT<31> ;
  wire \DSP_ALU.ALU_OUT<32> ;
  wire \DSP_ALU.ALU_OUT<33> ;
  wire \DSP_ALU.ALU_OUT<34> ;
  wire \DSP_ALU.ALU_OUT<35> ;
  wire \DSP_ALU.ALU_OUT<36> ;
  wire \DSP_ALU.ALU_OUT<37> ;
  wire \DSP_ALU.ALU_OUT<38> ;
  wire \DSP_ALU.ALU_OUT<39> ;
  wire \DSP_ALU.ALU_OUT<3> ;
  wire \DSP_ALU.ALU_OUT<40> ;
  wire \DSP_ALU.ALU_OUT<41> ;
  wire \DSP_ALU.ALU_OUT<42> ;
  wire \DSP_ALU.ALU_OUT<43> ;
  wire \DSP_ALU.ALU_OUT<44> ;
  wire \DSP_ALU.ALU_OUT<45> ;
  wire \DSP_ALU.ALU_OUT<46> ;
  wire \DSP_ALU.ALU_OUT<47> ;
  wire \DSP_ALU.ALU_OUT<4> ;
  wire \DSP_ALU.ALU_OUT<5> ;
  wire \DSP_ALU.ALU_OUT<6> ;
  wire \DSP_ALU.ALU_OUT<7> ;
  wire \DSP_ALU.ALU_OUT<8> ;
  wire \DSP_ALU.ALU_OUT<9> ;
  wire \DSP_ALU.COUT<0> ;
  wire \DSP_ALU.COUT<1> ;
  wire \DSP_ALU.COUT<2> ;
  wire \DSP_ALU.COUT<3> ;
  wire \DSP_ALU.MULTSIGN_ALU ;
  wire \DSP_ALU.XOR_MX<0> ;
  wire \DSP_ALU.XOR_MX<1> ;
  wire \DSP_ALU.XOR_MX<2> ;
  wire \DSP_ALU.XOR_MX<3> ;
  wire \DSP_ALU.XOR_MX<4> ;
  wire \DSP_ALU.XOR_MX<5> ;
  wire \DSP_ALU.XOR_MX<6> ;
  wire \DSP_ALU.XOR_MX<7> ;
  wire \DSP_A_B_DATA.A1_DATA<0> ;
  wire \DSP_A_B_DATA.A1_DATA<10> ;
  wire \DSP_A_B_DATA.A1_DATA<11> ;
  wire \DSP_A_B_DATA.A1_DATA<12> ;
  wire \DSP_A_B_DATA.A1_DATA<13> ;
  wire \DSP_A_B_DATA.A1_DATA<14> ;
  wire \DSP_A_B_DATA.A1_DATA<15> ;
  wire \DSP_A_B_DATA.A1_DATA<16> ;
  wire \DSP_A_B_DATA.A1_DATA<17> ;
  wire \DSP_A_B_DATA.A1_DATA<18> ;
  wire \DSP_A_B_DATA.A1_DATA<19> ;
  wire \DSP_A_B_DATA.A1_DATA<1> ;
  wire \DSP_A_B_DATA.A1_DATA<20> ;
  wire \DSP_A_B_DATA.A1_DATA<21> ;
  wire \DSP_A_B_DATA.A1_DATA<22> ;
  wire \DSP_A_B_DATA.A1_DATA<23> ;
  wire \DSP_A_B_DATA.A1_DATA<24> ;
  wire \DSP_A_B_DATA.A1_DATA<25> ;
  wire \DSP_A_B_DATA.A1_DATA<26> ;
  wire \DSP_A_B_DATA.A1_DATA<2> ;
  wire \DSP_A_B_DATA.A1_DATA<3> ;
  wire \DSP_A_B_DATA.A1_DATA<4> ;
  wire \DSP_A_B_DATA.A1_DATA<5> ;
  wire \DSP_A_B_DATA.A1_DATA<6> ;
  wire \DSP_A_B_DATA.A1_DATA<7> ;
  wire \DSP_A_B_DATA.A1_DATA<8> ;
  wire \DSP_A_B_DATA.A1_DATA<9> ;
  wire \DSP_A_B_DATA.A2_DATA<0> ;
  wire \DSP_A_B_DATA.A2_DATA<10> ;
  wire \DSP_A_B_DATA.A2_DATA<11> ;
  wire \DSP_A_B_DATA.A2_DATA<12> ;
  wire \DSP_A_B_DATA.A2_DATA<13> ;
  wire \DSP_A_B_DATA.A2_DATA<14> ;
  wire \DSP_A_B_DATA.A2_DATA<15> ;
  wire \DSP_A_B_DATA.A2_DATA<16> ;
  wire \DSP_A_B_DATA.A2_DATA<17> ;
  wire \DSP_A_B_DATA.A2_DATA<18> ;
  wire \DSP_A_B_DATA.A2_DATA<19> ;
  wire \DSP_A_B_DATA.A2_DATA<1> ;
  wire \DSP_A_B_DATA.A2_DATA<20> ;
  wire \DSP_A_B_DATA.A2_DATA<21> ;
  wire \DSP_A_B_DATA.A2_DATA<22> ;
  wire \DSP_A_B_DATA.A2_DATA<23> ;
  wire \DSP_A_B_DATA.A2_DATA<24> ;
  wire \DSP_A_B_DATA.A2_DATA<25> ;
  wire \DSP_A_B_DATA.A2_DATA<26> ;
  wire \DSP_A_B_DATA.A2_DATA<2> ;
  wire \DSP_A_B_DATA.A2_DATA<3> ;
  wire \DSP_A_B_DATA.A2_DATA<4> ;
  wire \DSP_A_B_DATA.A2_DATA<5> ;
  wire \DSP_A_B_DATA.A2_DATA<6> ;
  wire \DSP_A_B_DATA.A2_DATA<7> ;
  wire \DSP_A_B_DATA.A2_DATA<8> ;
  wire \DSP_A_B_DATA.A2_DATA<9> ;
  wire \DSP_A_B_DATA.A_ALU<0> ;
  wire \DSP_A_B_DATA.A_ALU<10> ;
  wire \DSP_A_B_DATA.A_ALU<11> ;
  wire \DSP_A_B_DATA.A_ALU<12> ;
  wire \DSP_A_B_DATA.A_ALU<13> ;
  wire \DSP_A_B_DATA.A_ALU<14> ;
  wire \DSP_A_B_DATA.A_ALU<15> ;
  wire \DSP_A_B_DATA.A_ALU<16> ;
  wire \DSP_A_B_DATA.A_ALU<17> ;
  wire \DSP_A_B_DATA.A_ALU<18> ;
  wire \DSP_A_B_DATA.A_ALU<19> ;
  wire \DSP_A_B_DATA.A_ALU<1> ;
  wire \DSP_A_B_DATA.A_ALU<20> ;
  wire \DSP_A_B_DATA.A_ALU<21> ;
  wire \DSP_A_B_DATA.A_ALU<22> ;
  wire \DSP_A_B_DATA.A_ALU<23> ;
  wire \DSP_A_B_DATA.A_ALU<24> ;
  wire \DSP_A_B_DATA.A_ALU<25> ;
  wire \DSP_A_B_DATA.A_ALU<26> ;
  wire \DSP_A_B_DATA.A_ALU<27> ;
  wire \DSP_A_B_DATA.A_ALU<28> ;
  wire \DSP_A_B_DATA.A_ALU<29> ;
  wire \DSP_A_B_DATA.A_ALU<2> ;
  wire \DSP_A_B_DATA.A_ALU<3> ;
  wire \DSP_A_B_DATA.A_ALU<4> ;
  wire \DSP_A_B_DATA.A_ALU<5> ;
  wire \DSP_A_B_DATA.A_ALU<6> ;
  wire \DSP_A_B_DATA.A_ALU<7> ;
  wire \DSP_A_B_DATA.A_ALU<8> ;
  wire \DSP_A_B_DATA.A_ALU<9> ;
  wire \DSP_A_B_DATA.B1_DATA<0> ;
  wire \DSP_A_B_DATA.B1_DATA<10> ;
  wire \DSP_A_B_DATA.B1_DATA<11> ;
  wire \DSP_A_B_DATA.B1_DATA<12> ;
  wire \DSP_A_B_DATA.B1_DATA<13> ;
  wire \DSP_A_B_DATA.B1_DATA<14> ;
  wire \DSP_A_B_DATA.B1_DATA<15> ;
  wire \DSP_A_B_DATA.B1_DATA<16> ;
  wire \DSP_A_B_DATA.B1_DATA<17> ;
  wire \DSP_A_B_DATA.B1_DATA<1> ;
  wire \DSP_A_B_DATA.B1_DATA<2> ;
  wire \DSP_A_B_DATA.B1_DATA<3> ;
  wire \DSP_A_B_DATA.B1_DATA<4> ;
  wire \DSP_A_B_DATA.B1_DATA<5> ;
  wire \DSP_A_B_DATA.B1_DATA<6> ;
  wire \DSP_A_B_DATA.B1_DATA<7> ;
  wire \DSP_A_B_DATA.B1_DATA<8> ;
  wire \DSP_A_B_DATA.B1_DATA<9> ;
  wire \DSP_A_B_DATA.B2_DATA<0> ;
  wire \DSP_A_B_DATA.B2_DATA<10> ;
  wire \DSP_A_B_DATA.B2_DATA<11> ;
  wire \DSP_A_B_DATA.B2_DATA<12> ;
  wire \DSP_A_B_DATA.B2_DATA<13> ;
  wire \DSP_A_B_DATA.B2_DATA<14> ;
  wire \DSP_A_B_DATA.B2_DATA<15> ;
  wire \DSP_A_B_DATA.B2_DATA<16> ;
  wire \DSP_A_B_DATA.B2_DATA<17> ;
  wire \DSP_A_B_DATA.B2_DATA<1> ;
  wire \DSP_A_B_DATA.B2_DATA<2> ;
  wire \DSP_A_B_DATA.B2_DATA<3> ;
  wire \DSP_A_B_DATA.B2_DATA<4> ;
  wire \DSP_A_B_DATA.B2_DATA<5> ;
  wire \DSP_A_B_DATA.B2_DATA<6> ;
  wire \DSP_A_B_DATA.B2_DATA<7> ;
  wire \DSP_A_B_DATA.B2_DATA<8> ;
  wire \DSP_A_B_DATA.B2_DATA<9> ;
  wire \DSP_A_B_DATA.B_ALU<0> ;
  wire \DSP_A_B_DATA.B_ALU<10> ;
  wire \DSP_A_B_DATA.B_ALU<11> ;
  wire \DSP_A_B_DATA.B_ALU<12> ;
  wire \DSP_A_B_DATA.B_ALU<13> ;
  wire \DSP_A_B_DATA.B_ALU<14> ;
  wire \DSP_A_B_DATA.B_ALU<15> ;
  wire \DSP_A_B_DATA.B_ALU<16> ;
  wire \DSP_A_B_DATA.B_ALU<17> ;
  wire \DSP_A_B_DATA.B_ALU<1> ;
  wire \DSP_A_B_DATA.B_ALU<2> ;
  wire \DSP_A_B_DATA.B_ALU<3> ;
  wire \DSP_A_B_DATA.B_ALU<4> ;
  wire \DSP_A_B_DATA.B_ALU<5> ;
  wire \DSP_A_B_DATA.B_ALU<6> ;
  wire \DSP_A_B_DATA.B_ALU<7> ;
  wire \DSP_A_B_DATA.B_ALU<8> ;
  wire \DSP_A_B_DATA.B_ALU<9> ;
  wire \DSP_C_DATA.C_DATA<0> ;
  wire \DSP_C_DATA.C_DATA<10> ;
  wire \DSP_C_DATA.C_DATA<11> ;
  wire \DSP_C_DATA.C_DATA<12> ;
  wire \DSP_C_DATA.C_DATA<13> ;
  wire \DSP_C_DATA.C_DATA<14> ;
  wire \DSP_C_DATA.C_DATA<15> ;
  wire \DSP_C_DATA.C_DATA<16> ;
  wire \DSP_C_DATA.C_DATA<17> ;
  wire \DSP_C_DATA.C_DATA<18> ;
  wire \DSP_C_DATA.C_DATA<19> ;
  wire \DSP_C_DATA.C_DATA<1> ;
  wire \DSP_C_DATA.C_DATA<20> ;
  wire \DSP_C_DATA.C_DATA<21> ;
  wire \DSP_C_DATA.C_DATA<22> ;
  wire \DSP_C_DATA.C_DATA<23> ;
  wire \DSP_C_DATA.C_DATA<24> ;
  wire \DSP_C_DATA.C_DATA<25> ;
  wire \DSP_C_DATA.C_DATA<26> ;
  wire \DSP_C_DATA.C_DATA<27> ;
  wire \DSP_C_DATA.C_DATA<28> ;
  wire \DSP_C_DATA.C_DATA<29> ;
  wire \DSP_C_DATA.C_DATA<2> ;
  wire \DSP_C_DATA.C_DATA<30> ;
  wire \DSP_C_DATA.C_DATA<31> ;
  wire \DSP_C_DATA.C_DATA<32> ;
  wire \DSP_C_DATA.C_DATA<33> ;
  wire \DSP_C_DATA.C_DATA<34> ;
  wire \DSP_C_DATA.C_DATA<35> ;
  wire \DSP_C_DATA.C_DATA<36> ;
  wire \DSP_C_DATA.C_DATA<37> ;
  wire \DSP_C_DATA.C_DATA<38> ;
  wire \DSP_C_DATA.C_DATA<39> ;
  wire \DSP_C_DATA.C_DATA<3> ;
  wire \DSP_C_DATA.C_DATA<40> ;
  wire \DSP_C_DATA.C_DATA<41> ;
  wire \DSP_C_DATA.C_DATA<42> ;
  wire \DSP_C_DATA.C_DATA<43> ;
  wire \DSP_C_DATA.C_DATA<44> ;
  wire \DSP_C_DATA.C_DATA<45> ;
  wire \DSP_C_DATA.C_DATA<46> ;
  wire \DSP_C_DATA.C_DATA<47> ;
  wire \DSP_C_DATA.C_DATA<4> ;
  wire \DSP_C_DATA.C_DATA<5> ;
  wire \DSP_C_DATA.C_DATA<6> ;
  wire \DSP_C_DATA.C_DATA<7> ;
  wire \DSP_C_DATA.C_DATA<8> ;
  wire \DSP_C_DATA.C_DATA<9> ;
  wire \DSP_MULTIPLIER.AMULT26 ;
  wire \DSP_MULTIPLIER.BMULT17 ;
  wire \DSP_MULTIPLIER.U<0> ;
  wire \DSP_MULTIPLIER.U<10> ;
  wire \DSP_MULTIPLIER.U<11> ;
  wire \DSP_MULTIPLIER.U<12> ;
  wire \DSP_MULTIPLIER.U<13> ;
  wire \DSP_MULTIPLIER.U<14> ;
  wire \DSP_MULTIPLIER.U<15> ;
  wire \DSP_MULTIPLIER.U<16> ;
  wire \DSP_MULTIPLIER.U<17> ;
  wire \DSP_MULTIPLIER.U<18> ;
  wire \DSP_MULTIPLIER.U<19> ;
  wire \DSP_MULTIPLIER.U<1> ;
  wire \DSP_MULTIPLIER.U<20> ;
  wire \DSP_MULTIPLIER.U<21> ;
  wire \DSP_MULTIPLIER.U<22> ;
  wire \DSP_MULTIPLIER.U<23> ;
  wire \DSP_MULTIPLIER.U<24> ;
  wire \DSP_MULTIPLIER.U<25> ;
  wire \DSP_MULTIPLIER.U<26> ;
  wire \DSP_MULTIPLIER.U<27> ;
  wire \DSP_MULTIPLIER.U<28> ;
  wire \DSP_MULTIPLIER.U<29> ;
  wire \DSP_MULTIPLIER.U<2> ;
  wire \DSP_MULTIPLIER.U<30> ;
  wire \DSP_MULTIPLIER.U<31> ;
  wire \DSP_MULTIPLIER.U<32> ;
  wire \DSP_MULTIPLIER.U<33> ;
  wire \DSP_MULTIPLIER.U<34> ;
  wire \DSP_MULTIPLIER.U<35> ;
  wire \DSP_MULTIPLIER.U<36> ;
  wire \DSP_MULTIPLIER.U<37> ;
  wire \DSP_MULTIPLIER.U<38> ;
  wire \DSP_MULTIPLIER.U<39> ;
  wire \DSP_MULTIPLIER.U<3> ;
  wire \DSP_MULTIPLIER.U<40> ;
  wire \DSP_MULTIPLIER.U<41> ;
  wire \DSP_MULTIPLIER.U<42> ;
  wire \DSP_MULTIPLIER.U<43> ;
  wire \DSP_MULTIPLIER.U<44> ;
  wire \DSP_MULTIPLIER.U<4> ;
  wire \DSP_MULTIPLIER.U<5> ;
  wire \DSP_MULTIPLIER.U<6> ;
  wire \DSP_MULTIPLIER.U<7> ;
  wire \DSP_MULTIPLIER.U<8> ;
  wire \DSP_MULTIPLIER.U<9> ;
  wire \DSP_MULTIPLIER.V<0> ;
  wire \DSP_MULTIPLIER.V<10> ;
  wire \DSP_MULTIPLIER.V<11> ;
  wire \DSP_MULTIPLIER.V<12> ;
  wire \DSP_MULTIPLIER.V<13> ;
  wire \DSP_MULTIPLIER.V<14> ;
  wire \DSP_MULTIPLIER.V<15> ;
  wire \DSP_MULTIPLIER.V<16> ;
  wire \DSP_MULTIPLIER.V<17> ;
  wire \DSP_MULTIPLIER.V<18> ;
  wire \DSP_MULTIPLIER.V<19> ;
  wire \DSP_MULTIPLIER.V<1> ;
  wire \DSP_MULTIPLIER.V<20> ;
  wire \DSP_MULTIPLIER.V<21> ;
  wire \DSP_MULTIPLIER.V<22> ;
  wire \DSP_MULTIPLIER.V<23> ;
  wire \DSP_MULTIPLIER.V<24> ;
  wire \DSP_MULTIPLIER.V<25> ;
  wire \DSP_MULTIPLIER.V<26> ;
  wire \DSP_MULTIPLIER.V<27> ;
  wire \DSP_MULTIPLIER.V<28> ;
  wire \DSP_MULTIPLIER.V<29> ;
  wire \DSP_MULTIPLIER.V<2> ;
  wire \DSP_MULTIPLIER.V<30> ;
  wire \DSP_MULTIPLIER.V<31> ;
  wire \DSP_MULTIPLIER.V<32> ;
  wire \DSP_MULTIPLIER.V<33> ;
  wire \DSP_MULTIPLIER.V<34> ;
  wire \DSP_MULTIPLIER.V<35> ;
  wire \DSP_MULTIPLIER.V<36> ;
  wire \DSP_MULTIPLIER.V<37> ;
  wire \DSP_MULTIPLIER.V<38> ;
  wire \DSP_MULTIPLIER.V<39> ;
  wire \DSP_MULTIPLIER.V<3> ;
  wire \DSP_MULTIPLIER.V<40> ;
  wire \DSP_MULTIPLIER.V<41> ;
  wire \DSP_MULTIPLIER.V<42> ;
  wire \DSP_MULTIPLIER.V<43> ;
  wire \DSP_MULTIPLIER.V<44> ;
  wire \DSP_MULTIPLIER.V<4> ;
  wire \DSP_MULTIPLIER.V<5> ;
  wire \DSP_MULTIPLIER.V<6> ;
  wire \DSP_MULTIPLIER.V<7> ;
  wire \DSP_MULTIPLIER.V<8> ;
  wire \DSP_MULTIPLIER.V<9> ;
  wire \DSP_M_DATA.U_DATA<0> ;
  wire \DSP_M_DATA.U_DATA<10> ;
  wire \DSP_M_DATA.U_DATA<11> ;
  wire \DSP_M_DATA.U_DATA<12> ;
  wire \DSP_M_DATA.U_DATA<13> ;
  wire \DSP_M_DATA.U_DATA<14> ;
  wire \DSP_M_DATA.U_DATA<15> ;
  wire \DSP_M_DATA.U_DATA<16> ;
  wire \DSP_M_DATA.U_DATA<17> ;
  wire \DSP_M_DATA.U_DATA<18> ;
  wire \DSP_M_DATA.U_DATA<19> ;
  wire \DSP_M_DATA.U_DATA<1> ;
  wire \DSP_M_DATA.U_DATA<20> ;
  wire \DSP_M_DATA.U_DATA<21> ;
  wire \DSP_M_DATA.U_DATA<22> ;
  wire \DSP_M_DATA.U_DATA<23> ;
  wire \DSP_M_DATA.U_DATA<24> ;
  wire \DSP_M_DATA.U_DATA<25> ;
  wire \DSP_M_DATA.U_DATA<26> ;
  wire \DSP_M_DATA.U_DATA<27> ;
  wire \DSP_M_DATA.U_DATA<28> ;
  wire \DSP_M_DATA.U_DATA<29> ;
  wire \DSP_M_DATA.U_DATA<2> ;
  wire \DSP_M_DATA.U_DATA<30> ;
  wire \DSP_M_DATA.U_DATA<31> ;
  wire \DSP_M_DATA.U_DATA<32> ;
  wire \DSP_M_DATA.U_DATA<33> ;
  wire \DSP_M_DATA.U_DATA<34> ;
  wire \DSP_M_DATA.U_DATA<35> ;
  wire \DSP_M_DATA.U_DATA<36> ;
  wire \DSP_M_DATA.U_DATA<37> ;
  wire \DSP_M_DATA.U_DATA<38> ;
  wire \DSP_M_DATA.U_DATA<39> ;
  wire \DSP_M_DATA.U_DATA<3> ;
  wire \DSP_M_DATA.U_DATA<40> ;
  wire \DSP_M_DATA.U_DATA<41> ;
  wire \DSP_M_DATA.U_DATA<42> ;
  wire \DSP_M_DATA.U_DATA<43> ;
  wire \DSP_M_DATA.U_DATA<44> ;
  wire \DSP_M_DATA.U_DATA<4> ;
  wire \DSP_M_DATA.U_DATA<5> ;
  wire \DSP_M_DATA.U_DATA<6> ;
  wire \DSP_M_DATA.U_DATA<7> ;
  wire \DSP_M_DATA.U_DATA<8> ;
  wire \DSP_M_DATA.U_DATA<9> ;
  wire \DSP_M_DATA.V_DATA<0> ;
  wire \DSP_M_DATA.V_DATA<10> ;
  wire \DSP_M_DATA.V_DATA<11> ;
  wire \DSP_M_DATA.V_DATA<12> ;
  wire \DSP_M_DATA.V_DATA<13> ;
  wire \DSP_M_DATA.V_DATA<14> ;
  wire \DSP_M_DATA.V_DATA<15> ;
  wire \DSP_M_DATA.V_DATA<16> ;
  wire \DSP_M_DATA.V_DATA<17> ;
  wire \DSP_M_DATA.V_DATA<18> ;
  wire \DSP_M_DATA.V_DATA<19> ;
  wire \DSP_M_DATA.V_DATA<1> ;
  wire \DSP_M_DATA.V_DATA<20> ;
  wire \DSP_M_DATA.V_DATA<21> ;
  wire \DSP_M_DATA.V_DATA<22> ;
  wire \DSP_M_DATA.V_DATA<23> ;
  wire \DSP_M_DATA.V_DATA<24> ;
  wire \DSP_M_DATA.V_DATA<25> ;
  wire \DSP_M_DATA.V_DATA<26> ;
  wire \DSP_M_DATA.V_DATA<27> ;
  wire \DSP_M_DATA.V_DATA<28> ;
  wire \DSP_M_DATA.V_DATA<29> ;
  wire \DSP_M_DATA.V_DATA<2> ;
  wire \DSP_M_DATA.V_DATA<30> ;
  wire \DSP_M_DATA.V_DATA<31> ;
  wire \DSP_M_DATA.V_DATA<32> ;
  wire \DSP_M_DATA.V_DATA<33> ;
  wire \DSP_M_DATA.V_DATA<34> ;
  wire \DSP_M_DATA.V_DATA<35> ;
  wire \DSP_M_DATA.V_DATA<36> ;
  wire \DSP_M_DATA.V_DATA<37> ;
  wire \DSP_M_DATA.V_DATA<38> ;
  wire \DSP_M_DATA.V_DATA<39> ;
  wire \DSP_M_DATA.V_DATA<3> ;
  wire \DSP_M_DATA.V_DATA<40> ;
  wire \DSP_M_DATA.V_DATA<41> ;
  wire \DSP_M_DATA.V_DATA<42> ;
  wire \DSP_M_DATA.V_DATA<43> ;
  wire \DSP_M_DATA.V_DATA<44> ;
  wire \DSP_M_DATA.V_DATA<4> ;
  wire \DSP_M_DATA.V_DATA<5> ;
  wire \DSP_M_DATA.V_DATA<6> ;
  wire \DSP_M_DATA.V_DATA<7> ;
  wire \DSP_M_DATA.V_DATA<8> ;
  wire \DSP_M_DATA.V_DATA<9> ;
  wire \DSP_OUTPUT.CCOUT_FB ;
  wire \DSP_OUTPUT.P_FDBK<0> ;
  wire \DSP_OUTPUT.P_FDBK<10> ;
  wire \DSP_OUTPUT.P_FDBK<11> ;
  wire \DSP_OUTPUT.P_FDBK<12> ;
  wire \DSP_OUTPUT.P_FDBK<13> ;
  wire \DSP_OUTPUT.P_FDBK<14> ;
  wire \DSP_OUTPUT.P_FDBK<15> ;
  wire \DSP_OUTPUT.P_FDBK<16> ;
  wire \DSP_OUTPUT.P_FDBK<17> ;
  wire \DSP_OUTPUT.P_FDBK<18> ;
  wire \DSP_OUTPUT.P_FDBK<19> ;
  wire \DSP_OUTPUT.P_FDBK<1> ;
  wire \DSP_OUTPUT.P_FDBK<20> ;
  wire \DSP_OUTPUT.P_FDBK<21> ;
  wire \DSP_OUTPUT.P_FDBK<22> ;
  wire \DSP_OUTPUT.P_FDBK<23> ;
  wire \DSP_OUTPUT.P_FDBK<24> ;
  wire \DSP_OUTPUT.P_FDBK<25> ;
  wire \DSP_OUTPUT.P_FDBK<26> ;
  wire \DSP_OUTPUT.P_FDBK<27> ;
  wire \DSP_OUTPUT.P_FDBK<28> ;
  wire \DSP_OUTPUT.P_FDBK<29> ;
  wire \DSP_OUTPUT.P_FDBK<2> ;
  wire \DSP_OUTPUT.P_FDBK<30> ;
  wire \DSP_OUTPUT.P_FDBK<31> ;
  wire \DSP_OUTPUT.P_FDBK<32> ;
  wire \DSP_OUTPUT.P_FDBK<33> ;
  wire \DSP_OUTPUT.P_FDBK<34> ;
  wire \DSP_OUTPUT.P_FDBK<35> ;
  wire \DSP_OUTPUT.P_FDBK<36> ;
  wire \DSP_OUTPUT.P_FDBK<37> ;
  wire \DSP_OUTPUT.P_FDBK<38> ;
  wire \DSP_OUTPUT.P_FDBK<39> ;
  wire \DSP_OUTPUT.P_FDBK<3> ;
  wire \DSP_OUTPUT.P_FDBK<40> ;
  wire \DSP_OUTPUT.P_FDBK<41> ;
  wire \DSP_OUTPUT.P_FDBK<42> ;
  wire \DSP_OUTPUT.P_FDBK<43> ;
  wire \DSP_OUTPUT.P_FDBK<44> ;
  wire \DSP_OUTPUT.P_FDBK<45> ;
  wire \DSP_OUTPUT.P_FDBK<46> ;
  wire \DSP_OUTPUT.P_FDBK<47> ;
  wire \DSP_OUTPUT.P_FDBK<4> ;
  wire \DSP_OUTPUT.P_FDBK<5> ;
  wire \DSP_OUTPUT.P_FDBK<6> ;
  wire \DSP_OUTPUT.P_FDBK<7> ;
  wire \DSP_OUTPUT.P_FDBK<8> ;
  wire \DSP_OUTPUT.P_FDBK<9> ;
  wire \DSP_OUTPUT.P_FDBK_47 ;
  wire \DSP_PREADD.AD<0> ;
  wire \DSP_PREADD.AD<10> ;
  wire \DSP_PREADD.AD<11> ;
  wire \DSP_PREADD.AD<12> ;
  wire \DSP_PREADD.AD<13> ;
  wire \DSP_PREADD.AD<14> ;
  wire \DSP_PREADD.AD<15> ;
  wire \DSP_PREADD.AD<16> ;
  wire \DSP_PREADD.AD<17> ;
  wire \DSP_PREADD.AD<18> ;
  wire \DSP_PREADD.AD<19> ;
  wire \DSP_PREADD.AD<1> ;
  wire \DSP_PREADD.AD<20> ;
  wire \DSP_PREADD.AD<21> ;
  wire \DSP_PREADD.AD<22> ;
  wire \DSP_PREADD.AD<23> ;
  wire \DSP_PREADD.AD<24> ;
  wire \DSP_PREADD.AD<25> ;
  wire \DSP_PREADD.AD<26> ;
  wire \DSP_PREADD.AD<2> ;
  wire \DSP_PREADD.AD<3> ;
  wire \DSP_PREADD.AD<4> ;
  wire \DSP_PREADD.AD<5> ;
  wire \DSP_PREADD.AD<6> ;
  wire \DSP_PREADD.AD<7> ;
  wire \DSP_PREADD.AD<8> ;
  wire \DSP_PREADD.AD<9> ;
  wire \DSP_PREADD_DATA.A2A1<0> ;
  wire \DSP_PREADD_DATA.A2A1<10> ;
  wire \DSP_PREADD_DATA.A2A1<11> ;
  wire \DSP_PREADD_DATA.A2A1<12> ;
  wire \DSP_PREADD_DATA.A2A1<13> ;
  wire \DSP_PREADD_DATA.A2A1<14> ;
  wire \DSP_PREADD_DATA.A2A1<15> ;
  wire \DSP_PREADD_DATA.A2A1<16> ;
  wire \DSP_PREADD_DATA.A2A1<17> ;
  wire \DSP_PREADD_DATA.A2A1<18> ;
  wire \DSP_PREADD_DATA.A2A1<19> ;
  wire \DSP_PREADD_DATA.A2A1<1> ;
  wire \DSP_PREADD_DATA.A2A1<20> ;
  wire \DSP_PREADD_DATA.A2A1<21> ;
  wire \DSP_PREADD_DATA.A2A1<22> ;
  wire \DSP_PREADD_DATA.A2A1<23> ;
  wire \DSP_PREADD_DATA.A2A1<24> ;
  wire \DSP_PREADD_DATA.A2A1<25> ;
  wire \DSP_PREADD_DATA.A2A1<26> ;
  wire \DSP_PREADD_DATA.A2A1<2> ;
  wire \DSP_PREADD_DATA.A2A1<3> ;
  wire \DSP_PREADD_DATA.A2A1<4> ;
  wire \DSP_PREADD_DATA.A2A1<5> ;
  wire \DSP_PREADD_DATA.A2A1<6> ;
  wire \DSP_PREADD_DATA.A2A1<7> ;
  wire \DSP_PREADD_DATA.A2A1<8> ;
  wire \DSP_PREADD_DATA.A2A1<9> ;
  wire \DSP_PREADD_DATA.ADDSUB ;
  wire \DSP_PREADD_DATA.AD_DATA<0> ;
  wire \DSP_PREADD_DATA.AD_DATA<10> ;
  wire \DSP_PREADD_DATA.AD_DATA<11> ;
  wire \DSP_PREADD_DATA.AD_DATA<12> ;
  wire \DSP_PREADD_DATA.AD_DATA<13> ;
  wire \DSP_PREADD_DATA.AD_DATA<14> ;
  wire \DSP_PREADD_DATA.AD_DATA<15> ;
  wire \DSP_PREADD_DATA.AD_DATA<16> ;
  wire \DSP_PREADD_DATA.AD_DATA<17> ;
  wire \DSP_PREADD_DATA.AD_DATA<18> ;
  wire \DSP_PREADD_DATA.AD_DATA<19> ;
  wire \DSP_PREADD_DATA.AD_DATA<1> ;
  wire \DSP_PREADD_DATA.AD_DATA<20> ;
  wire \DSP_PREADD_DATA.AD_DATA<21> ;
  wire \DSP_PREADD_DATA.AD_DATA<22> ;
  wire \DSP_PREADD_DATA.AD_DATA<23> ;
  wire \DSP_PREADD_DATA.AD_DATA<24> ;
  wire \DSP_PREADD_DATA.AD_DATA<25> ;
  wire \DSP_PREADD_DATA.AD_DATA<26> ;
  wire \DSP_PREADD_DATA.AD_DATA<2> ;
  wire \DSP_PREADD_DATA.AD_DATA<3> ;
  wire \DSP_PREADD_DATA.AD_DATA<4> ;
  wire \DSP_PREADD_DATA.AD_DATA<5> ;
  wire \DSP_PREADD_DATA.AD_DATA<6> ;
  wire \DSP_PREADD_DATA.AD_DATA<7> ;
  wire \DSP_PREADD_DATA.AD_DATA<8> ;
  wire \DSP_PREADD_DATA.AD_DATA<9> ;
  wire \DSP_PREADD_DATA.B2B1<0> ;
  wire \DSP_PREADD_DATA.B2B1<10> ;
  wire \DSP_PREADD_DATA.B2B1<11> ;
  wire \DSP_PREADD_DATA.B2B1<12> ;
  wire \DSP_PREADD_DATA.B2B1<13> ;
  wire \DSP_PREADD_DATA.B2B1<14> ;
  wire \DSP_PREADD_DATA.B2B1<15> ;
  wire \DSP_PREADD_DATA.B2B1<16> ;
  wire \DSP_PREADD_DATA.B2B1<17> ;
  wire \DSP_PREADD_DATA.B2B1<1> ;
  wire \DSP_PREADD_DATA.B2B1<2> ;
  wire \DSP_PREADD_DATA.B2B1<3> ;
  wire \DSP_PREADD_DATA.B2B1<4> ;
  wire \DSP_PREADD_DATA.B2B1<5> ;
  wire \DSP_PREADD_DATA.B2B1<6> ;
  wire \DSP_PREADD_DATA.B2B1<7> ;
  wire \DSP_PREADD_DATA.B2B1<8> ;
  wire \DSP_PREADD_DATA.B2B1<9> ;
  wire \DSP_PREADD_DATA.D_DATA<0> ;
  wire \DSP_PREADD_DATA.D_DATA<10> ;
  wire \DSP_PREADD_DATA.D_DATA<11> ;
  wire \DSP_PREADD_DATA.D_DATA<12> ;
  wire \DSP_PREADD_DATA.D_DATA<13> ;
  wire \DSP_PREADD_DATA.D_DATA<14> ;
  wire \DSP_PREADD_DATA.D_DATA<15> ;
  wire \DSP_PREADD_DATA.D_DATA<16> ;
  wire \DSP_PREADD_DATA.D_DATA<17> ;
  wire \DSP_PREADD_DATA.D_DATA<18> ;
  wire \DSP_PREADD_DATA.D_DATA<19> ;
  wire \DSP_PREADD_DATA.D_DATA<1> ;
  wire \DSP_PREADD_DATA.D_DATA<20> ;
  wire \DSP_PREADD_DATA.D_DATA<21> ;
  wire \DSP_PREADD_DATA.D_DATA<22> ;
  wire \DSP_PREADD_DATA.D_DATA<23> ;
  wire \DSP_PREADD_DATA.D_DATA<24> ;
  wire \DSP_PREADD_DATA.D_DATA<25> ;
  wire \DSP_PREADD_DATA.D_DATA<26> ;
  wire \DSP_PREADD_DATA.D_DATA<2> ;
  wire \DSP_PREADD_DATA.D_DATA<3> ;
  wire \DSP_PREADD_DATA.D_DATA<4> ;
  wire \DSP_PREADD_DATA.D_DATA<5> ;
  wire \DSP_PREADD_DATA.D_DATA<6> ;
  wire \DSP_PREADD_DATA.D_DATA<7> ;
  wire \DSP_PREADD_DATA.D_DATA<8> ;
  wire \DSP_PREADD_DATA.D_DATA<9> ;
  wire \DSP_PREADD_DATA.INMODE_2 ;
  wire \DSP_PREADD_DATA.PREADD_AB<0> ;
  wire \DSP_PREADD_DATA.PREADD_AB<10> ;
  wire \DSP_PREADD_DATA.PREADD_AB<11> ;
  wire \DSP_PREADD_DATA.PREADD_AB<12> ;
  wire \DSP_PREADD_DATA.PREADD_AB<13> ;
  wire \DSP_PREADD_DATA.PREADD_AB<14> ;
  wire \DSP_PREADD_DATA.PREADD_AB<15> ;
  wire \DSP_PREADD_DATA.PREADD_AB<16> ;
  wire \DSP_PREADD_DATA.PREADD_AB<17> ;
  wire \DSP_PREADD_DATA.PREADD_AB<18> ;
  wire \DSP_PREADD_DATA.PREADD_AB<19> ;
  wire \DSP_PREADD_DATA.PREADD_AB<1> ;
  wire \DSP_PREADD_DATA.PREADD_AB<20> ;
  wire \DSP_PREADD_DATA.PREADD_AB<21> ;
  wire \DSP_PREADD_DATA.PREADD_AB<22> ;
  wire \DSP_PREADD_DATA.PREADD_AB<23> ;
  wire \DSP_PREADD_DATA.PREADD_AB<24> ;
  wire \DSP_PREADD_DATA.PREADD_AB<25> ;
  wire \DSP_PREADD_DATA.PREADD_AB<26> ;
  wire \DSP_PREADD_DATA.PREADD_AB<2> ;
  wire \DSP_PREADD_DATA.PREADD_AB<3> ;
  wire \DSP_PREADD_DATA.PREADD_AB<4> ;
  wire \DSP_PREADD_DATA.PREADD_AB<5> ;
  wire \DSP_PREADD_DATA.PREADD_AB<6> ;
  wire \DSP_PREADD_DATA.PREADD_AB<7> ;
  wire \DSP_PREADD_DATA.PREADD_AB<8> ;
  wire \DSP_PREADD_DATA.PREADD_AB<9> ;
  wire \D[0] ;
  wire \D[10] ;
  wire \D[11] ;
  wire \D[12] ;
  wire \D[13] ;
  wire \D[14] ;
  wire \D[15] ;
  wire \D[16] ;
  wire \D[17] ;
  wire \D[18] ;
  wire \D[19] ;
  wire \D[1] ;
  wire \D[20] ;
  wire \D[21] ;
  wire \D[22] ;
  wire \D[23] ;
  wire \D[24] ;
  wire \D[25] ;
  wire \D[26] ;
  wire \D[2] ;
  wire \D[3] ;
  wire \D[4] ;
  wire \D[5] ;
  wire \D[6] ;
  wire \D[7] ;
  wire \D[8] ;
  wire \D[9] ;
  wire \INMODE[0] ;
  wire \INMODE[1] ;
  wire \INMODE[2] ;
  wire \INMODE[3] ;
  wire \INMODE[4] ;
  wire MULTSIGNIN;
  wire MULTSIGNOUT;
  wire \OPMODE[0] ;
  wire \OPMODE[1] ;
  wire \OPMODE[2] ;
  wire \OPMODE[3] ;
  wire \OPMODE[4] ;
  wire \OPMODE[5] ;
  wire \OPMODE[6] ;
  wire \OPMODE[7] ;
  wire \OPMODE[8] ;
  wire OVERFLOW;
  wire PATTERNBDETECT;
  wire PATTERNDETECT;
  wire \PCIN[0] ;
  wire \PCIN[10] ;
  wire \PCIN[11] ;
  wire \PCIN[12] ;
  wire \PCIN[13] ;
  wire \PCIN[14] ;
  wire \PCIN[15] ;
  wire \PCIN[16] ;
  wire \PCIN[17] ;
  wire \PCIN[18] ;
  wire \PCIN[19] ;
  wire \PCIN[1] ;
  wire \PCIN[20] ;
  wire \PCIN[21] ;
  wire \PCIN[22] ;
  wire \PCIN[23] ;
  wire \PCIN[24] ;
  wire \PCIN[25] ;
  wire \PCIN[26] ;
  wire \PCIN[27] ;
  wire \PCIN[28] ;
  wire \PCIN[29] ;
  wire \PCIN[2] ;
  wire \PCIN[30] ;
  wire \PCIN[31] ;
  wire \PCIN[32] ;
  wire \PCIN[33] ;
  wire \PCIN[34] ;
  wire \PCIN[35] ;
  wire \PCIN[36] ;
  wire \PCIN[37] ;
  wire \PCIN[38] ;
  wire \PCIN[39] ;
  wire \PCIN[3] ;
  wire \PCIN[40] ;
  wire \PCIN[41] ;
  wire \PCIN[42] ;
  wire \PCIN[43] ;
  wire \PCIN[44] ;
  wire \PCIN[45] ;
  wire \PCIN[46] ;
  wire \PCIN[47] ;
  wire \PCIN[4] ;
  wire \PCIN[5] ;
  wire \PCIN[6] ;
  wire \PCIN[7] ;
  wire \PCIN[8] ;
  wire \PCIN[9] ;
  wire \PCOUT[0] ;
  wire \PCOUT[10] ;
  wire \PCOUT[11] ;
  wire \PCOUT[12] ;
  wire \PCOUT[13] ;
  wire \PCOUT[14] ;
  wire \PCOUT[15] ;
  wire \PCOUT[16] ;
  wire \PCOUT[17] ;
  wire \PCOUT[18] ;
  wire \PCOUT[19] ;
  wire \PCOUT[1] ;
  wire \PCOUT[20] ;
  wire \PCOUT[21] ;
  wire \PCOUT[22] ;
  wire \PCOUT[23] ;
  wire \PCOUT[24] ;
  wire \PCOUT[25] ;
  wire \PCOUT[26] ;
  wire \PCOUT[27] ;
  wire \PCOUT[28] ;
  wire \PCOUT[29] ;
  wire \PCOUT[2] ;
  wire \PCOUT[30] ;
  wire \PCOUT[31] ;
  wire \PCOUT[32] ;
  wire \PCOUT[33] ;
  wire \PCOUT[34] ;
  wire \PCOUT[35] ;
  wire \PCOUT[36] ;
  wire \PCOUT[37] ;
  wire \PCOUT[38] ;
  wire \PCOUT[39] ;
  wire \PCOUT[3] ;
  wire \PCOUT[40] ;
  wire \PCOUT[41] ;
  wire \PCOUT[42] ;
  wire \PCOUT[43] ;
  wire \PCOUT[44] ;
  wire \PCOUT[45] ;
  wire \PCOUT[46] ;
  wire \PCOUT[47] ;
  wire \PCOUT[4] ;
  wire \PCOUT[5] ;
  wire \PCOUT[6] ;
  wire \PCOUT[7] ;
  wire \PCOUT[8] ;
  wire \PCOUT[9] ;
  wire \P[0] ;
  wire \P[10] ;
  wire \P[11] ;
  wire \P[12] ;
  wire \P[13] ;
  wire \P[14] ;
  wire \P[15] ;
  wire \P[16] ;
  wire \P[17] ;
  wire \P[18] ;
  wire \P[19] ;
  wire \P[1] ;
  wire \P[20] ;
  wire \P[21] ;
  wire \P[22] ;
  wire \P[23] ;
  wire \P[24] ;
  wire \P[25] ;
  wire \P[26] ;
  wire \P[27] ;
  wire \P[28] ;
  wire \P[29] ;
  wire \P[2] ;
  wire \P[30] ;
  wire \P[31] ;
  wire \P[32] ;
  wire \P[33] ;
  wire \P[34] ;
  wire \P[35] ;
  wire \P[36] ;
  wire \P[37] ;
  wire \P[38] ;
  wire \P[39] ;
  wire \P[3] ;
  wire \P[40] ;
  wire \P[41] ;
  wire \P[42] ;
  wire \P[43] ;
  wire \P[44] ;
  wire \P[45] ;
  wire \P[46] ;
  wire \P[47] ;
  wire \P[4] ;
  wire \P[5] ;
  wire \P[6] ;
  wire \P[7] ;
  wire \P[8] ;
  wire \P[9] ;
  wire RSTA;
  wire RSTALLCARRYIN;
  wire RSTALUMODE;
  wire RSTB;
  wire RSTC;
  wire RSTCTRL;
  wire RSTD;
  wire RSTINMODE;
  wire RSTM;
  wire RSTP;
  wire UNDERFLOW;
  wire \XOROUT[0] ;
  wire \XOROUT[1] ;
  wire \XOROUT[2] ;
  wire \XOROUT[3] ;
  wire \XOROUT[4] ;
  wire \XOROUT[5] ;
  wire \XOROUT[6] ;
  wire \XOROUT[7] ;

  assign \ACIN[0]  = ACIN[0];
  assign \ACIN[10]  = ACIN[10];
  assign \ACIN[11]  = ACIN[11];
  assign \ACIN[12]  = ACIN[12];
  assign \ACIN[13]  = ACIN[13];
  assign \ACIN[14]  = ACIN[14];
  assign \ACIN[15]  = ACIN[15];
  assign \ACIN[16]  = ACIN[16];
  assign \ACIN[17]  = ACIN[17];
  assign \ACIN[18]  = ACIN[18];
  assign \ACIN[19]  = ACIN[19];
  assign \ACIN[1]  = ACIN[1];
  assign \ACIN[20]  = ACIN[20];
  assign \ACIN[21]  = ACIN[21];
  assign \ACIN[22]  = ACIN[22];
  assign \ACIN[23]  = ACIN[23];
  assign \ACIN[24]  = ACIN[24];
  assign \ACIN[25]  = ACIN[25];
  assign \ACIN[26]  = ACIN[26];
  assign \ACIN[27]  = ACIN[27];
  assign \ACIN[28]  = ACIN[28];
  assign \ACIN[29]  = ACIN[29];
  assign \ACIN[2]  = ACIN[2];
  assign \ACIN[3]  = ACIN[3];
  assign \ACIN[4]  = ACIN[4];
  assign \ACIN[5]  = ACIN[5];
  assign \ACIN[6]  = ACIN[6];
  assign \ACIN[7]  = ACIN[7];
  assign \ACIN[8]  = ACIN[8];
  assign \ACIN[9]  = ACIN[9];
  assign ACOUT[29] = \ACOUT[29] ;
  assign ACOUT[28] = \ACOUT[28] ;
  assign ACOUT[27] = \ACOUT[27] ;
  assign ACOUT[26] = \ACOUT[26] ;
  assign ACOUT[25] = \ACOUT[25] ;
  assign ACOUT[24] = \ACOUT[24] ;
  assign ACOUT[23] = \ACOUT[23] ;
  assign ACOUT[22] = \ACOUT[22] ;
  assign ACOUT[21] = \ACOUT[21] ;
  assign ACOUT[20] = \ACOUT[20] ;
  assign ACOUT[19] = \ACOUT[19] ;
  assign ACOUT[18] = \ACOUT[18] ;
  assign ACOUT[17] = \ACOUT[17] ;
  assign ACOUT[16] = \ACOUT[16] ;
  assign ACOUT[15] = \ACOUT[15] ;
  assign ACOUT[14] = \ACOUT[14] ;
  assign ACOUT[13] = \ACOUT[13] ;
  assign ACOUT[12] = \ACOUT[12] ;
  assign ACOUT[11] = \ACOUT[11] ;
  assign ACOUT[10] = \ACOUT[10] ;
  assign ACOUT[9] = \ACOUT[9] ;
  assign ACOUT[8] = \ACOUT[8] ;
  assign ACOUT[7] = \ACOUT[7] ;
  assign ACOUT[6] = \ACOUT[6] ;
  assign ACOUT[5] = \ACOUT[5] ;
  assign ACOUT[4] = \ACOUT[4] ;
  assign ACOUT[3] = \ACOUT[3] ;
  assign ACOUT[2] = \ACOUT[2] ;
  assign ACOUT[1] = \ACOUT[1] ;
  assign ACOUT[0] = \ACOUT[0] ;
  assign \ALUMODE[0]  = ALUMODE[0];
  assign \ALUMODE[1]  = ALUMODE[1];
  assign \ALUMODE[2]  = ALUMODE[2];
  assign \ALUMODE[3]  = ALUMODE[3];
  assign \A[0]  = A[0];
  assign \A[10]  = A[10];
  assign \A[11]  = A[11];
  assign \A[12]  = A[12];
  assign \A[13]  = A[13];
  assign \A[14]  = A[14];
  assign \A[15]  = A[15];
  assign \A[16]  = A[16];
  assign \A[17]  = A[17];
  assign \A[18]  = A[18];
  assign \A[19]  = A[19];
  assign \A[1]  = A[1];
  assign \A[20]  = A[20];
  assign \A[21]  = A[21];
  assign \A[22]  = A[22];
  assign \A[23]  = A[23];
  assign \A[24]  = A[24];
  assign \A[25]  = A[25];
  assign \A[26]  = A[26];
  assign \A[27]  = A[27];
  assign \A[28]  = A[28];
  assign \A[29]  = A[29];
  assign \A[2]  = A[2];
  assign \A[3]  = A[3];
  assign \A[4]  = A[4];
  assign \A[5]  = A[5];
  assign \A[6]  = A[6];
  assign \A[7]  = A[7];
  assign \A[8]  = A[8];
  assign \A[9]  = A[9];
  assign \BCIN[0]  = BCIN[0];
  assign \BCIN[10]  = BCIN[10];
  assign \BCIN[11]  = BCIN[11];
  assign \BCIN[12]  = BCIN[12];
  assign \BCIN[13]  = BCIN[13];
  assign \BCIN[14]  = BCIN[14];
  assign \BCIN[15]  = BCIN[15];
  assign \BCIN[16]  = BCIN[16];
  assign \BCIN[17]  = BCIN[17];
  assign \BCIN[1]  = BCIN[1];
  assign \BCIN[2]  = BCIN[2];
  assign \BCIN[3]  = BCIN[3];
  assign \BCIN[4]  = BCIN[4];
  assign \BCIN[5]  = BCIN[5];
  assign \BCIN[6]  = BCIN[6];
  assign \BCIN[7]  = BCIN[7];
  assign \BCIN[8]  = BCIN[8];
  assign \BCIN[9]  = BCIN[9];
  assign BCOUT[17] = \BCOUT[17] ;
  assign BCOUT[16] = \BCOUT[16] ;
  assign BCOUT[15] = \BCOUT[15] ;
  assign BCOUT[14] = \BCOUT[14] ;
  assign BCOUT[13] = \BCOUT[13] ;
  assign BCOUT[12] = \BCOUT[12] ;
  assign BCOUT[11] = \BCOUT[11] ;
  assign BCOUT[10] = \BCOUT[10] ;
  assign BCOUT[9] = \BCOUT[9] ;
  assign BCOUT[8] = \BCOUT[8] ;
  assign BCOUT[7] = \BCOUT[7] ;
  assign BCOUT[6] = \BCOUT[6] ;
  assign BCOUT[5] = \BCOUT[5] ;
  assign BCOUT[4] = \BCOUT[4] ;
  assign BCOUT[3] = \BCOUT[3] ;
  assign BCOUT[2] = \BCOUT[2] ;
  assign BCOUT[1] = \BCOUT[1] ;
  assign BCOUT[0] = \BCOUT[0] ;
  assign \B[0]  = B[0];
  assign \B[10]  = B[10];
  assign \B[11]  = B[11];
  assign \B[12]  = B[12];
  assign \B[13]  = B[13];
  assign \B[14]  = B[14];
  assign \B[15]  = B[15];
  assign \B[16]  = B[16];
  assign \B[17]  = B[17];
  assign \B[1]  = B[1];
  assign \B[2]  = B[2];
  assign \B[3]  = B[3];
  assign \B[4]  = B[4];
  assign \B[5]  = B[5];
  assign \B[6]  = B[6];
  assign \B[7]  = B[7];
  assign \B[8]  = B[8];
  assign \B[9]  = B[9];
  assign \CARRYINSEL[0]  = CARRYINSEL[0];
  assign \CARRYINSEL[1]  = CARRYINSEL[1];
  assign \CARRYINSEL[2]  = CARRYINSEL[2];
  assign CARRYOUT[3] = \CARRYOUT[3] ;
  assign CARRYOUT[2] = \CARRYOUT[2] ;
  assign CARRYOUT[1] = \CARRYOUT[1] ;
  assign CARRYOUT[0] = \CARRYOUT[0] ;
  assign \C[0]  = C[0];
  assign \C[10]  = C[10];
  assign \C[11]  = C[11];
  assign \C[12]  = C[12];
  assign \C[13]  = C[13];
  assign \C[14]  = C[14];
  assign \C[15]  = C[15];
  assign \C[16]  = C[16];
  assign \C[17]  = C[17];
  assign \C[18]  = C[18];
  assign \C[19]  = C[19];
  assign \C[1]  = C[1];
  assign \C[20]  = C[20];
  assign \C[21]  = C[21];
  assign \C[22]  = C[22];
  assign \C[23]  = C[23];
  assign \C[24]  = C[24];
  assign \C[25]  = C[25];
  assign \C[26]  = C[26];
  assign \C[27]  = C[27];
  assign \C[28]  = C[28];
  assign \C[29]  = C[29];
  assign \C[2]  = C[2];
  assign \C[30]  = C[30];
  assign \C[31]  = C[31];
  assign \C[32]  = C[32];
  assign \C[33]  = C[33];
  assign \C[34]  = C[34];
  assign \C[35]  = C[35];
  assign \C[36]  = C[36];
  assign \C[37]  = C[37];
  assign \C[38]  = C[38];
  assign \C[39]  = C[39];
  assign \C[3]  = C[3];
  assign \C[40]  = C[40];
  assign \C[41]  = C[41];
  assign \C[42]  = C[42];
  assign \C[43]  = C[43];
  assign \C[44]  = C[44];
  assign \C[45]  = C[45];
  assign \C[46]  = C[46];
  assign \C[47]  = C[47];
  assign \C[4]  = C[4];
  assign \C[5]  = C[5];
  assign \C[6]  = C[6];
  assign \C[7]  = C[7];
  assign \C[8]  = C[8];
  assign \C[9]  = C[9];
  assign \D[0]  = D[0];
  assign \D[10]  = D[10];
  assign \D[11]  = D[11];
  assign \D[12]  = D[12];
  assign \D[13]  = D[13];
  assign \D[14]  = D[14];
  assign \D[15]  = D[15];
  assign \D[16]  = D[16];
  assign \D[17]  = D[17];
  assign \D[18]  = D[18];
  assign \D[19]  = D[19];
  assign \D[1]  = D[1];
  assign \D[20]  = D[20];
  assign \D[21]  = D[21];
  assign \D[22]  = D[22];
  assign \D[23]  = D[23];
  assign \D[24]  = D[24];
  assign \D[25]  = D[25];
  assign \D[26]  = D[26];
  assign \D[2]  = D[2];
  assign \D[3]  = D[3];
  assign \D[4]  = D[4];
  assign \D[5]  = D[5];
  assign \D[6]  = D[6];
  assign \D[7]  = D[7];
  assign \D[8]  = D[8];
  assign \D[9]  = D[9];
  assign \INMODE[0]  = INMODE[0];
  assign \INMODE[1]  = INMODE[1];
  assign \INMODE[2]  = INMODE[2];
  assign \INMODE[3]  = INMODE[3];
  assign \INMODE[4]  = INMODE[4];
  assign \OPMODE[0]  = OPMODE[0];
  assign \OPMODE[1]  = OPMODE[1];
  assign \OPMODE[2]  = OPMODE[2];
  assign \OPMODE[3]  = OPMODE[3];
  assign \OPMODE[4]  = OPMODE[4];
  assign \OPMODE[5]  = OPMODE[5];
  assign \OPMODE[6]  = OPMODE[6];
  assign \OPMODE[7]  = OPMODE[7];
  assign \OPMODE[8]  = OPMODE[8];
  assign P[47] = \P[47] ;
  assign P[46] = \P[46] ;
  assign P[45] = \P[45] ;
  assign P[44] = \P[44] ;
  assign P[43] = \P[43] ;
  assign P[42] = \P[42] ;
  assign P[41] = \P[41] ;
  assign P[40] = \P[40] ;
  assign P[39] = \P[39] ;
  assign P[38] = \P[38] ;
  assign P[37] = \P[37] ;
  assign P[36] = \P[36] ;
  assign P[35] = \P[35] ;
  assign P[34] = \P[34] ;
  assign P[33] = \P[33] ;
  assign P[32] = \P[32] ;
  assign P[31] = \P[31] ;
  assign P[30] = \P[30] ;
  assign P[29] = \P[29] ;
  assign P[28] = \P[28] ;
  assign P[27] = \P[27] ;
  assign P[26] = \P[26] ;
  assign P[25] = \P[25] ;
  assign P[24] = \P[24] ;
  assign P[23] = \P[23] ;
  assign P[22] = \P[22] ;
  assign P[21] = \P[21] ;
  assign P[20] = \P[20] ;
  assign P[19] = \P[19] ;
  assign P[18] = \P[18] ;
  assign P[17] = \P[17] ;
  assign P[16] = \P[16] ;
  assign P[15] = \P[15] ;
  assign P[14] = \P[14] ;
  assign P[13] = \P[13] ;
  assign P[12] = \P[12] ;
  assign P[11] = \P[11] ;
  assign P[10] = \P[10] ;
  assign P[9] = \P[9] ;
  assign P[8] = \P[8] ;
  assign P[7] = \P[7] ;
  assign P[6] = \P[6] ;
  assign P[5] = \P[5] ;
  assign P[4] = \P[4] ;
  assign P[3] = \P[3] ;
  assign P[2] = \P[2] ;
  assign P[1] = \P[1] ;
  assign P[0] = \P[0] ;
  assign \PCIN[0]  = PCIN[0];
  assign \PCIN[10]  = PCIN[10];
  assign \PCIN[11]  = PCIN[11];
  assign \PCIN[12]  = PCIN[12];
  assign \PCIN[13]  = PCIN[13];
  assign \PCIN[14]  = PCIN[14];
  assign \PCIN[15]  = PCIN[15];
  assign \PCIN[16]  = PCIN[16];
  assign \PCIN[17]  = PCIN[17];
  assign \PCIN[18]  = PCIN[18];
  assign \PCIN[19]  = PCIN[19];
  assign \PCIN[1]  = PCIN[1];
  assign \PCIN[20]  = PCIN[20];
  assign \PCIN[21]  = PCIN[21];
  assign \PCIN[22]  = PCIN[22];
  assign \PCIN[23]  = PCIN[23];
  assign \PCIN[24]  = PCIN[24];
  assign \PCIN[25]  = PCIN[25];
  assign \PCIN[26]  = PCIN[26];
  assign \PCIN[27]  = PCIN[27];
  assign \PCIN[28]  = PCIN[28];
  assign \PCIN[29]  = PCIN[29];
  assign \PCIN[2]  = PCIN[2];
  assign \PCIN[30]  = PCIN[30];
  assign \PCIN[31]  = PCIN[31];
  assign \PCIN[32]  = PCIN[32];
  assign \PCIN[33]  = PCIN[33];
  assign \PCIN[34]  = PCIN[34];
  assign \PCIN[35]  = PCIN[35];
  assign \PCIN[36]  = PCIN[36];
  assign \PCIN[37]  = PCIN[37];
  assign \PCIN[38]  = PCIN[38];
  assign \PCIN[39]  = PCIN[39];
  assign \PCIN[3]  = PCIN[3];
  assign \PCIN[40]  = PCIN[40];
  assign \PCIN[41]  = PCIN[41];
  assign \PCIN[42]  = PCIN[42];
  assign \PCIN[43]  = PCIN[43];
  assign \PCIN[44]  = PCIN[44];
  assign \PCIN[45]  = PCIN[45];
  assign \PCIN[46]  = PCIN[46];
  assign \PCIN[47]  = PCIN[47];
  assign \PCIN[4]  = PCIN[4];
  assign \PCIN[5]  = PCIN[5];
  assign \PCIN[6]  = PCIN[6];
  assign \PCIN[7]  = PCIN[7];
  assign \PCIN[8]  = PCIN[8];
  assign \PCIN[9]  = PCIN[9];
  assign PCOUT[47] = \PCOUT[47] ;
  assign PCOUT[46] = \PCOUT[46] ;
  assign PCOUT[45] = \PCOUT[45] ;
  assign PCOUT[44] = \PCOUT[44] ;
  assign PCOUT[43] = \PCOUT[43] ;
  assign PCOUT[42] = \PCOUT[42] ;
  assign PCOUT[41] = \PCOUT[41] ;
  assign PCOUT[40] = \PCOUT[40] ;
  assign PCOUT[39] = \PCOUT[39] ;
  assign PCOUT[38] = \PCOUT[38] ;
  assign PCOUT[37] = \PCOUT[37] ;
  assign PCOUT[36] = \PCOUT[36] ;
  assign PCOUT[35] = \PCOUT[35] ;
  assign PCOUT[34] = \PCOUT[34] ;
  assign PCOUT[33] = \PCOUT[33] ;
  assign PCOUT[32] = \PCOUT[32] ;
  assign PCOUT[31] = \PCOUT[31] ;
  assign PCOUT[30] = \PCOUT[30] ;
  assign PCOUT[29] = \PCOUT[29] ;
  assign PCOUT[28] = \PCOUT[28] ;
  assign PCOUT[27] = \PCOUT[27] ;
  assign PCOUT[26] = \PCOUT[26] ;
  assign PCOUT[25] = \PCOUT[25] ;
  assign PCOUT[24] = \PCOUT[24] ;
  assign PCOUT[23] = \PCOUT[23] ;
  assign PCOUT[22] = \PCOUT[22] ;
  assign PCOUT[21] = \PCOUT[21] ;
  assign PCOUT[20] = \PCOUT[20] ;
  assign PCOUT[19] = \PCOUT[19] ;
  assign PCOUT[18] = \PCOUT[18] ;
  assign PCOUT[17] = \PCOUT[17] ;
  assign PCOUT[16] = \PCOUT[16] ;
  assign PCOUT[15] = \PCOUT[15] ;
  assign PCOUT[14] = \PCOUT[14] ;
  assign PCOUT[13] = \PCOUT[13] ;
  assign PCOUT[12] = \PCOUT[12] ;
  assign PCOUT[11] = \PCOUT[11] ;
  assign PCOUT[10] = \PCOUT[10] ;
  assign PCOUT[9] = \PCOUT[9] ;
  assign PCOUT[8] = \PCOUT[8] ;
  assign PCOUT[7] = \PCOUT[7] ;
  assign PCOUT[6] = \PCOUT[6] ;
  assign PCOUT[5] = \PCOUT[5] ;
  assign PCOUT[4] = \PCOUT[4] ;
  assign PCOUT[3] = \PCOUT[3] ;
  assign PCOUT[2] = \PCOUT[2] ;
  assign PCOUT[1] = \PCOUT[1] ;
  assign PCOUT[0] = \PCOUT[0] ;
  assign XOROUT[7] = \XOROUT[7] ;
  assign XOROUT[6] = \XOROUT[6] ;
  assign XOROUT[5] = \XOROUT[5] ;
  assign XOROUT[4] = \XOROUT[4] ;
  assign XOROUT[3] = \XOROUT[3] ;
  assign XOROUT[2] = \XOROUT[2] ;
  assign XOROUT[1] = \XOROUT[1] ;
  assign XOROUT[0] = \XOROUT[0] ;
  DSP_ALU #(
    .ALUMODEREG(0),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_OPMODE_INVERTED(9'b000000000),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .MREG(0),
    .OPMODEREG(0),
    .RND(48'h000000000000),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")) 
    DSP_ALU_INST
       (.ALUMODE({\ALUMODE[3] ,\ALUMODE[2] ,\ALUMODE[1] ,\ALUMODE[0] }),
        .ALUMODE10(\DSP_ALU.ALUMODE10 ),
        .ALU_OUT({\DSP_ALU.ALU_OUT<47> ,\DSP_ALU.ALU_OUT<46> ,\DSP_ALU.ALU_OUT<45> ,\DSP_ALU.ALU_OUT<44> ,\DSP_ALU.ALU_OUT<43> ,\DSP_ALU.ALU_OUT<42> ,\DSP_ALU.ALU_OUT<41> ,\DSP_ALU.ALU_OUT<40> ,\DSP_ALU.ALU_OUT<39> ,\DSP_ALU.ALU_OUT<38> ,\DSP_ALU.ALU_OUT<37> ,\DSP_ALU.ALU_OUT<36> ,\DSP_ALU.ALU_OUT<35> ,\DSP_ALU.ALU_OUT<34> ,\DSP_ALU.ALU_OUT<33> ,\DSP_ALU.ALU_OUT<32> ,\DSP_ALU.ALU_OUT<31> ,\DSP_ALU.ALU_OUT<30> ,\DSP_ALU.ALU_OUT<29> ,\DSP_ALU.ALU_OUT<28> ,\DSP_ALU.ALU_OUT<27> ,\DSP_ALU.ALU_OUT<26> ,\DSP_ALU.ALU_OUT<25> ,\DSP_ALU.ALU_OUT<24> ,\DSP_ALU.ALU_OUT<23> ,\DSP_ALU.ALU_OUT<22> ,\DSP_ALU.ALU_OUT<21> ,\DSP_ALU.ALU_OUT<20> ,\DSP_ALU.ALU_OUT<19> ,\DSP_ALU.ALU_OUT<18> ,\DSP_ALU.ALU_OUT<17> ,\DSP_ALU.ALU_OUT<16> ,\DSP_ALU.ALU_OUT<15> ,\DSP_ALU.ALU_OUT<14> ,\DSP_ALU.ALU_OUT<13> ,\DSP_ALU.ALU_OUT<12> ,\DSP_ALU.ALU_OUT<11> ,\DSP_ALU.ALU_OUT<10> ,\DSP_ALU.ALU_OUT<9> ,\DSP_ALU.ALU_OUT<8> ,\DSP_ALU.ALU_OUT<7> ,\DSP_ALU.ALU_OUT<6> ,\DSP_ALU.ALU_OUT<5> ,\DSP_ALU.ALU_OUT<4> ,\DSP_ALU.ALU_OUT<3> ,\DSP_ALU.ALU_OUT<2> ,\DSP_ALU.ALU_OUT<1> ,\DSP_ALU.ALU_OUT<0> }),
        .AMULT26(\DSP_MULTIPLIER.AMULT26 ),
        .A_ALU({\DSP_A_B_DATA.A_ALU<29> ,\DSP_A_B_DATA.A_ALU<28> ,\DSP_A_B_DATA.A_ALU<27> ,\DSP_A_B_DATA.A_ALU<26> ,\DSP_A_B_DATA.A_ALU<25> ,\DSP_A_B_DATA.A_ALU<24> ,\DSP_A_B_DATA.A_ALU<23> ,\DSP_A_B_DATA.A_ALU<22> ,\DSP_A_B_DATA.A_ALU<21> ,\DSP_A_B_DATA.A_ALU<20> ,\DSP_A_B_DATA.A_ALU<19> ,\DSP_A_B_DATA.A_ALU<18> ,\DSP_A_B_DATA.A_ALU<17> ,\DSP_A_B_DATA.A_ALU<16> ,\DSP_A_B_DATA.A_ALU<15> ,\DSP_A_B_DATA.A_ALU<14> ,\DSP_A_B_DATA.A_ALU<13> ,\DSP_A_B_DATA.A_ALU<12> ,\DSP_A_B_DATA.A_ALU<11> ,\DSP_A_B_DATA.A_ALU<10> ,\DSP_A_B_DATA.A_ALU<9> ,\DSP_A_B_DATA.A_ALU<8> ,\DSP_A_B_DATA.A_ALU<7> ,\DSP_A_B_DATA.A_ALU<6> ,\DSP_A_B_DATA.A_ALU<5> ,\DSP_A_B_DATA.A_ALU<4> ,\DSP_A_B_DATA.A_ALU<3> ,\DSP_A_B_DATA.A_ALU<2> ,\DSP_A_B_DATA.A_ALU<1> ,\DSP_A_B_DATA.A_ALU<0> }),
        .BMULT17(\DSP_MULTIPLIER.BMULT17 ),
        .B_ALU({\DSP_A_B_DATA.B_ALU<17> ,\DSP_A_B_DATA.B_ALU<16> ,\DSP_A_B_DATA.B_ALU<15> ,\DSP_A_B_DATA.B_ALU<14> ,\DSP_A_B_DATA.B_ALU<13> ,\DSP_A_B_DATA.B_ALU<12> ,\DSP_A_B_DATA.B_ALU<11> ,\DSP_A_B_DATA.B_ALU<10> ,\DSP_A_B_DATA.B_ALU<9> ,\DSP_A_B_DATA.B_ALU<8> ,\DSP_A_B_DATA.B_ALU<7> ,\DSP_A_B_DATA.B_ALU<6> ,\DSP_A_B_DATA.B_ALU<5> ,\DSP_A_B_DATA.B_ALU<4> ,\DSP_A_B_DATA.B_ALU<3> ,\DSP_A_B_DATA.B_ALU<2> ,\DSP_A_B_DATA.B_ALU<1> ,\DSP_A_B_DATA.B_ALU<0> }),
        .CARRYCASCIN(CARRYCASCIN),
        .CARRYIN(CARRYIN),
        .CARRYINSEL({\CARRYINSEL[2] ,\CARRYINSEL[1] ,\CARRYINSEL[0] }),
        .CCOUT(\DSP_OUTPUT.CCOUT_FB ),
        .CEALUMODE(CEALUMODE),
        .CECARRYIN(CECARRYIN),
        .CECTRL(CECTRL),
        .CEM(CEM),
        .CLK(CLK),
        .COUT({\DSP_ALU.COUT<3> ,\DSP_ALU.COUT<2> ,\DSP_ALU.COUT<1> ,\DSP_ALU.COUT<0> }),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .MULTSIGNIN(MULTSIGNIN),
        .MULTSIGN_ALU(\DSP_ALU.MULTSIGN_ALU ),
        .OPMODE({\OPMODE[8] ,\OPMODE[7] ,\OPMODE[6] ,\OPMODE[5] ,\OPMODE[4] ,\OPMODE[3] ,\OPMODE[2] ,\OPMODE[1] ,\OPMODE[0] }),
        .PCIN({\PCIN[47] ,\PCIN[46] ,\PCIN[45] ,\PCIN[44] ,\PCIN[43] ,\PCIN[42] ,\PCIN[41] ,\PCIN[40] ,\PCIN[39] ,\PCIN[38] ,\PCIN[37] ,\PCIN[36] ,\PCIN[35] ,\PCIN[34] ,\PCIN[33] ,\PCIN[32] ,\PCIN[31] ,\PCIN[30] ,\PCIN[29] ,\PCIN[28] ,\PCIN[27] ,\PCIN[26] ,\PCIN[25] ,\PCIN[24] ,\PCIN[23] ,\PCIN[22] ,\PCIN[21] ,\PCIN[20] ,\PCIN[19] ,\PCIN[18] ,\PCIN[17] ,\PCIN[16] ,\PCIN[15] ,\PCIN[14] ,\PCIN[13] ,\PCIN[12] ,\PCIN[11] ,\PCIN[10] ,\PCIN[9] ,\PCIN[8] ,\PCIN[7] ,\PCIN[6] ,\PCIN[5] ,\PCIN[4] ,\PCIN[3] ,\PCIN[2] ,\PCIN[1] ,\PCIN[0] }),
        .P_FDBK({\DSP_OUTPUT.P_FDBK<47> ,\DSP_OUTPUT.P_FDBK<46> ,\DSP_OUTPUT.P_FDBK<45> ,\DSP_OUTPUT.P_FDBK<44> ,\DSP_OUTPUT.P_FDBK<43> ,\DSP_OUTPUT.P_FDBK<42> ,\DSP_OUTPUT.P_FDBK<41> ,\DSP_OUTPUT.P_FDBK<40> ,\DSP_OUTPUT.P_FDBK<39> ,\DSP_OUTPUT.P_FDBK<38> ,\DSP_OUTPUT.P_FDBK<37> ,\DSP_OUTPUT.P_FDBK<36> ,\DSP_OUTPUT.P_FDBK<35> ,\DSP_OUTPUT.P_FDBK<34> ,\DSP_OUTPUT.P_FDBK<33> ,\DSP_OUTPUT.P_FDBK<32> ,\DSP_OUTPUT.P_FDBK<31> ,\DSP_OUTPUT.P_FDBK<30> ,\DSP_OUTPUT.P_FDBK<29> ,\DSP_OUTPUT.P_FDBK<28> ,\DSP_OUTPUT.P_FDBK<27> ,\DSP_OUTPUT.P_FDBK<26> ,\DSP_OUTPUT.P_FDBK<25> ,\DSP_OUTPUT.P_FDBK<24> ,\DSP_OUTPUT.P_FDBK<23> ,\DSP_OUTPUT.P_FDBK<22> ,\DSP_OUTPUT.P_FDBK<21> ,\DSP_OUTPUT.P_FDBK<20> ,\DSP_OUTPUT.P_FDBK<19> ,\DSP_OUTPUT.P_FDBK<18> ,\DSP_OUTPUT.P_FDBK<17> ,\DSP_OUTPUT.P_FDBK<16> ,\DSP_OUTPUT.P_FDBK<15> ,\DSP_OUTPUT.P_FDBK<14> ,\DSP_OUTPUT.P_FDBK<13> ,\DSP_OUTPUT.P_FDBK<12> ,\DSP_OUTPUT.P_FDBK<11> ,\DSP_OUTPUT.P_FDBK<10> ,\DSP_OUTPUT.P_FDBK<9> ,\DSP_OUTPUT.P_FDBK<8> ,\DSP_OUTPUT.P_FDBK<7> ,\DSP_OUTPUT.P_FDBK<6> ,\DSP_OUTPUT.P_FDBK<5> ,\DSP_OUTPUT.P_FDBK<4> ,\DSP_OUTPUT.P_FDBK<3> ,\DSP_OUTPUT.P_FDBK<2> ,\DSP_OUTPUT.P_FDBK<1> ,\DSP_OUTPUT.P_FDBK<0> }),
        .P_FDBK_47(\DSP_OUTPUT.P_FDBK_47 ),
        .RSTALLCARRYIN(RSTALLCARRYIN),
        .RSTALUMODE(RSTALUMODE),
        .RSTCTRL(RSTCTRL),
        .U_DATA({\DSP_M_DATA.U_DATA<44> ,\DSP_M_DATA.U_DATA<43> ,\DSP_M_DATA.U_DATA<42> ,\DSP_M_DATA.U_DATA<41> ,\DSP_M_DATA.U_DATA<40> ,\DSP_M_DATA.U_DATA<39> ,\DSP_M_DATA.U_DATA<38> ,\DSP_M_DATA.U_DATA<37> ,\DSP_M_DATA.U_DATA<36> ,\DSP_M_DATA.U_DATA<35> ,\DSP_M_DATA.U_DATA<34> ,\DSP_M_DATA.U_DATA<33> ,\DSP_M_DATA.U_DATA<32> ,\DSP_M_DATA.U_DATA<31> ,\DSP_M_DATA.U_DATA<30> ,\DSP_M_DATA.U_DATA<29> ,\DSP_M_DATA.U_DATA<28> ,\DSP_M_DATA.U_DATA<27> ,\DSP_M_DATA.U_DATA<26> ,\DSP_M_DATA.U_DATA<25> ,\DSP_M_DATA.U_DATA<24> ,\DSP_M_DATA.U_DATA<23> ,\DSP_M_DATA.U_DATA<22> ,\DSP_M_DATA.U_DATA<21> ,\DSP_M_DATA.U_DATA<20> ,\DSP_M_DATA.U_DATA<19> ,\DSP_M_DATA.U_DATA<18> ,\DSP_M_DATA.U_DATA<17> ,\DSP_M_DATA.U_DATA<16> ,\DSP_M_DATA.U_DATA<15> ,\DSP_M_DATA.U_DATA<14> ,\DSP_M_DATA.U_DATA<13> ,\DSP_M_DATA.U_DATA<12> ,\DSP_M_DATA.U_DATA<11> ,\DSP_M_DATA.U_DATA<10> ,\DSP_M_DATA.U_DATA<9> ,\DSP_M_DATA.U_DATA<8> ,\DSP_M_DATA.U_DATA<7> ,\DSP_M_DATA.U_DATA<6> ,\DSP_M_DATA.U_DATA<5> ,\DSP_M_DATA.U_DATA<4> ,\DSP_M_DATA.U_DATA<3> ,\DSP_M_DATA.U_DATA<2> ,\DSP_M_DATA.U_DATA<1> ,\DSP_M_DATA.U_DATA<0> }),
        .V_DATA({\DSP_M_DATA.V_DATA<44> ,\DSP_M_DATA.V_DATA<43> ,\DSP_M_DATA.V_DATA<42> ,\DSP_M_DATA.V_DATA<41> ,\DSP_M_DATA.V_DATA<40> ,\DSP_M_DATA.V_DATA<39> ,\DSP_M_DATA.V_DATA<38> ,\DSP_M_DATA.V_DATA<37> ,\DSP_M_DATA.V_DATA<36> ,\DSP_M_DATA.V_DATA<35> ,\DSP_M_DATA.V_DATA<34> ,\DSP_M_DATA.V_DATA<33> ,\DSP_M_DATA.V_DATA<32> ,\DSP_M_DATA.V_DATA<31> ,\DSP_M_DATA.V_DATA<30> ,\DSP_M_DATA.V_DATA<29> ,\DSP_M_DATA.V_DATA<28> ,\DSP_M_DATA.V_DATA<27> ,\DSP_M_DATA.V_DATA<26> ,\DSP_M_DATA.V_DATA<25> ,\DSP_M_DATA.V_DATA<24> ,\DSP_M_DATA.V_DATA<23> ,\DSP_M_DATA.V_DATA<22> ,\DSP_M_DATA.V_DATA<21> ,\DSP_M_DATA.V_DATA<20> ,\DSP_M_DATA.V_DATA<19> ,\DSP_M_DATA.V_DATA<18> ,\DSP_M_DATA.V_DATA<17> ,\DSP_M_DATA.V_DATA<16> ,\DSP_M_DATA.V_DATA<15> ,\DSP_M_DATA.V_DATA<14> ,\DSP_M_DATA.V_DATA<13> ,\DSP_M_DATA.V_DATA<12> ,\DSP_M_DATA.V_DATA<11> ,\DSP_M_DATA.V_DATA<10> ,\DSP_M_DATA.V_DATA<9> ,\DSP_M_DATA.V_DATA<8> ,\DSP_M_DATA.V_DATA<7> ,\DSP_M_DATA.V_DATA<6> ,\DSP_M_DATA.V_DATA<5> ,\DSP_M_DATA.V_DATA<4> ,\DSP_M_DATA.V_DATA<3> ,\DSP_M_DATA.V_DATA<2> ,\DSP_M_DATA.V_DATA<1> ,\DSP_M_DATA.V_DATA<0> }),
        .XOR_MX({\DSP_ALU.XOR_MX<7> ,\DSP_ALU.XOR_MX<6> ,\DSP_ALU.XOR_MX<5> ,\DSP_ALU.XOR_MX<4> ,\DSP_ALU.XOR_MX<3> ,\DSP_ALU.XOR_MX<2> ,\DSP_ALU.XOR_MX<1> ,\DSP_ALU.XOR_MX<0> }));
  DSP_A_B_DATA #(
    .ACASCREG(0),
    .AREG(0),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0)) 
    DSP_A_B_DATA_INST
       (.A({\A[29] ,\A[28] ,\A[27] ,\A[26] ,\A[25] ,\A[24] ,\A[23] ,\A[22] ,\A[21] ,\A[20] ,\A[19] ,\A[18] ,\A[17] ,\A[16] ,\A[15] ,\A[14] ,\A[13] ,\A[12] ,\A[11] ,\A[10] ,\A[9] ,\A[8] ,\A[7] ,\A[6] ,\A[5] ,\A[4] ,\A[3] ,\A[2] ,\A[1] ,\A[0] }),
        .A1_DATA({\DSP_A_B_DATA.A1_DATA<26> ,\DSP_A_B_DATA.A1_DATA<25> ,\DSP_A_B_DATA.A1_DATA<24> ,\DSP_A_B_DATA.A1_DATA<23> ,\DSP_A_B_DATA.A1_DATA<22> ,\DSP_A_B_DATA.A1_DATA<21> ,\DSP_A_B_DATA.A1_DATA<20> ,\DSP_A_B_DATA.A1_DATA<19> ,\DSP_A_B_DATA.A1_DATA<18> ,\DSP_A_B_DATA.A1_DATA<17> ,\DSP_A_B_DATA.A1_DATA<16> ,\DSP_A_B_DATA.A1_DATA<15> ,\DSP_A_B_DATA.A1_DATA<14> ,\DSP_A_B_DATA.A1_DATA<13> ,\DSP_A_B_DATA.A1_DATA<12> ,\DSP_A_B_DATA.A1_DATA<11> ,\DSP_A_B_DATA.A1_DATA<10> ,\DSP_A_B_DATA.A1_DATA<9> ,\DSP_A_B_DATA.A1_DATA<8> ,\DSP_A_B_DATA.A1_DATA<7> ,\DSP_A_B_DATA.A1_DATA<6> ,\DSP_A_B_DATA.A1_DATA<5> ,\DSP_A_B_DATA.A1_DATA<4> ,\DSP_A_B_DATA.A1_DATA<3> ,\DSP_A_B_DATA.A1_DATA<2> ,\DSP_A_B_DATA.A1_DATA<1> ,\DSP_A_B_DATA.A1_DATA<0> }),
        .A2_DATA({\DSP_A_B_DATA.A2_DATA<26> ,\DSP_A_B_DATA.A2_DATA<25> ,\DSP_A_B_DATA.A2_DATA<24> ,\DSP_A_B_DATA.A2_DATA<23> ,\DSP_A_B_DATA.A2_DATA<22> ,\DSP_A_B_DATA.A2_DATA<21> ,\DSP_A_B_DATA.A2_DATA<20> ,\DSP_A_B_DATA.A2_DATA<19> ,\DSP_A_B_DATA.A2_DATA<18> ,\DSP_A_B_DATA.A2_DATA<17> ,\DSP_A_B_DATA.A2_DATA<16> ,\DSP_A_B_DATA.A2_DATA<15> ,\DSP_A_B_DATA.A2_DATA<14> ,\DSP_A_B_DATA.A2_DATA<13> ,\DSP_A_B_DATA.A2_DATA<12> ,\DSP_A_B_DATA.A2_DATA<11> ,\DSP_A_B_DATA.A2_DATA<10> ,\DSP_A_B_DATA.A2_DATA<9> ,\DSP_A_B_DATA.A2_DATA<8> ,\DSP_A_B_DATA.A2_DATA<7> ,\DSP_A_B_DATA.A2_DATA<6> ,\DSP_A_B_DATA.A2_DATA<5> ,\DSP_A_B_DATA.A2_DATA<4> ,\DSP_A_B_DATA.A2_DATA<3> ,\DSP_A_B_DATA.A2_DATA<2> ,\DSP_A_B_DATA.A2_DATA<1> ,\DSP_A_B_DATA.A2_DATA<0> }),
        .ACIN({\ACIN[29] ,\ACIN[28] ,\ACIN[27] ,\ACIN[26] ,\ACIN[25] ,\ACIN[24] ,\ACIN[23] ,\ACIN[22] ,\ACIN[21] ,\ACIN[20] ,\ACIN[19] ,\ACIN[18] ,\ACIN[17] ,\ACIN[16] ,\ACIN[15] ,\ACIN[14] ,\ACIN[13] ,\ACIN[12] ,\ACIN[11] ,\ACIN[10] ,\ACIN[9] ,\ACIN[8] ,\ACIN[7] ,\ACIN[6] ,\ACIN[5] ,\ACIN[4] ,\ACIN[3] ,\ACIN[2] ,\ACIN[1] ,\ACIN[0] }),
        .ACOUT({\ACOUT[29] ,\ACOUT[28] ,\ACOUT[27] ,\ACOUT[26] ,\ACOUT[25] ,\ACOUT[24] ,\ACOUT[23] ,\ACOUT[22] ,\ACOUT[21] ,\ACOUT[20] ,\ACOUT[19] ,\ACOUT[18] ,\ACOUT[17] ,\ACOUT[16] ,\ACOUT[15] ,\ACOUT[14] ,\ACOUT[13] ,\ACOUT[12] ,\ACOUT[11] ,\ACOUT[10] ,\ACOUT[9] ,\ACOUT[8] ,\ACOUT[7] ,\ACOUT[6] ,\ACOUT[5] ,\ACOUT[4] ,\ACOUT[3] ,\ACOUT[2] ,\ACOUT[1] ,\ACOUT[0] }),
        .A_ALU({\DSP_A_B_DATA.A_ALU<29> ,\DSP_A_B_DATA.A_ALU<28> ,\DSP_A_B_DATA.A_ALU<27> ,\DSP_A_B_DATA.A_ALU<26> ,\DSP_A_B_DATA.A_ALU<25> ,\DSP_A_B_DATA.A_ALU<24> ,\DSP_A_B_DATA.A_ALU<23> ,\DSP_A_B_DATA.A_ALU<22> ,\DSP_A_B_DATA.A_ALU<21> ,\DSP_A_B_DATA.A_ALU<20> ,\DSP_A_B_DATA.A_ALU<19> ,\DSP_A_B_DATA.A_ALU<18> ,\DSP_A_B_DATA.A_ALU<17> ,\DSP_A_B_DATA.A_ALU<16> ,\DSP_A_B_DATA.A_ALU<15> ,\DSP_A_B_DATA.A_ALU<14> ,\DSP_A_B_DATA.A_ALU<13> ,\DSP_A_B_DATA.A_ALU<12> ,\DSP_A_B_DATA.A_ALU<11> ,\DSP_A_B_DATA.A_ALU<10> ,\DSP_A_B_DATA.A_ALU<9> ,\DSP_A_B_DATA.A_ALU<8> ,\DSP_A_B_DATA.A_ALU<7> ,\DSP_A_B_DATA.A_ALU<6> ,\DSP_A_B_DATA.A_ALU<5> ,\DSP_A_B_DATA.A_ALU<4> ,\DSP_A_B_DATA.A_ALU<3> ,\DSP_A_B_DATA.A_ALU<2> ,\DSP_A_B_DATA.A_ALU<1> ,\DSP_A_B_DATA.A_ALU<0> }),
        .B({\B[17] ,\B[16] ,\B[15] ,\B[14] ,\B[13] ,\B[12] ,\B[11] ,\B[10] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,\B[0] }),
        .B1_DATA({\DSP_A_B_DATA.B1_DATA<17> ,\DSP_A_B_DATA.B1_DATA<16> ,\DSP_A_B_DATA.B1_DATA<15> ,\DSP_A_B_DATA.B1_DATA<14> ,\DSP_A_B_DATA.B1_DATA<13> ,\DSP_A_B_DATA.B1_DATA<12> ,\DSP_A_B_DATA.B1_DATA<11> ,\DSP_A_B_DATA.B1_DATA<10> ,\DSP_A_B_DATA.B1_DATA<9> ,\DSP_A_B_DATA.B1_DATA<8> ,\DSP_A_B_DATA.B1_DATA<7> ,\DSP_A_B_DATA.B1_DATA<6> ,\DSP_A_B_DATA.B1_DATA<5> ,\DSP_A_B_DATA.B1_DATA<4> ,\DSP_A_B_DATA.B1_DATA<3> ,\DSP_A_B_DATA.B1_DATA<2> ,\DSP_A_B_DATA.B1_DATA<1> ,\DSP_A_B_DATA.B1_DATA<0> }),
        .B2_DATA({\DSP_A_B_DATA.B2_DATA<17> ,\DSP_A_B_DATA.B2_DATA<16> ,\DSP_A_B_DATA.B2_DATA<15> ,\DSP_A_B_DATA.B2_DATA<14> ,\DSP_A_B_DATA.B2_DATA<13> ,\DSP_A_B_DATA.B2_DATA<12> ,\DSP_A_B_DATA.B2_DATA<11> ,\DSP_A_B_DATA.B2_DATA<10> ,\DSP_A_B_DATA.B2_DATA<9> ,\DSP_A_B_DATA.B2_DATA<8> ,\DSP_A_B_DATA.B2_DATA<7> ,\DSP_A_B_DATA.B2_DATA<6> ,\DSP_A_B_DATA.B2_DATA<5> ,\DSP_A_B_DATA.B2_DATA<4> ,\DSP_A_B_DATA.B2_DATA<3> ,\DSP_A_B_DATA.B2_DATA<2> ,\DSP_A_B_DATA.B2_DATA<1> ,\DSP_A_B_DATA.B2_DATA<0> }),
        .BCIN({\BCIN[17] ,\BCIN[16] ,\BCIN[15] ,\BCIN[14] ,\BCIN[13] ,\BCIN[12] ,\BCIN[11] ,\BCIN[10] ,\BCIN[9] ,\BCIN[8] ,\BCIN[7] ,\BCIN[6] ,\BCIN[5] ,\BCIN[4] ,\BCIN[3] ,\BCIN[2] ,\BCIN[1] ,\BCIN[0] }),
        .BCOUT({\BCOUT[17] ,\BCOUT[16] ,\BCOUT[15] ,\BCOUT[14] ,\BCOUT[13] ,\BCOUT[12] ,\BCOUT[11] ,\BCOUT[10] ,\BCOUT[9] ,\BCOUT[8] ,\BCOUT[7] ,\BCOUT[6] ,\BCOUT[5] ,\BCOUT[4] ,\BCOUT[3] ,\BCOUT[2] ,\BCOUT[1] ,\BCOUT[0] }),
        .B_ALU({\DSP_A_B_DATA.B_ALU<17> ,\DSP_A_B_DATA.B_ALU<16> ,\DSP_A_B_DATA.B_ALU<15> ,\DSP_A_B_DATA.B_ALU<14> ,\DSP_A_B_DATA.B_ALU<13> ,\DSP_A_B_DATA.B_ALU<12> ,\DSP_A_B_DATA.B_ALU<11> ,\DSP_A_B_DATA.B_ALU<10> ,\DSP_A_B_DATA.B_ALU<9> ,\DSP_A_B_DATA.B_ALU<8> ,\DSP_A_B_DATA.B_ALU<7> ,\DSP_A_B_DATA.B_ALU<6> ,\DSP_A_B_DATA.B_ALU<5> ,\DSP_A_B_DATA.B_ALU<4> ,\DSP_A_B_DATA.B_ALU<3> ,\DSP_A_B_DATA.B_ALU<2> ,\DSP_A_B_DATA.B_ALU<1> ,\DSP_A_B_DATA.B_ALU<0> }),
        .CEA1(CEA1),
        .CEA2(CEA2),
        .CEB1(CEB1),
        .CEB2(CEB2),
        .CLK(CLK),
        .RSTA(RSTA),
        .RSTB(RSTB));
  DSP_C_DATA #(
    .CREG(0),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0)) 
    DSP_C_DATA_INST
       (.C({\C[47] ,\C[46] ,\C[45] ,\C[44] ,\C[43] ,\C[42] ,\C[41] ,\C[40] ,\C[39] ,\C[38] ,\C[37] ,\C[36] ,\C[35] ,\C[34] ,\C[33] ,\C[32] ,\C[31] ,\C[30] ,\C[29] ,\C[28] ,\C[27] ,\C[26] ,\C[25] ,\C[24] ,\C[23] ,\C[22] ,\C[21] ,\C[20] ,\C[19] ,\C[18] ,\C[17] ,\C[16] ,\C[15] ,\C[14] ,\C[13] ,\C[12] ,\C[11] ,\C[10] ,\C[9] ,\C[8] ,\C[7] ,\C[6] ,\C[5] ,\C[4] ,\C[3] ,\C[2] ,\C[1] ,\C[0] }),
        .CEC(CEC),
        .CLK(CLK),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .RSTC(RSTC));
  DSP_MULTIPLIER #(
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .USE_MULT("MULTIPLY")) 
    DSP_MULTIPLIER_INST
       (.A2A1({\DSP_PREADD_DATA.A2A1<26> ,\DSP_PREADD_DATA.A2A1<25> ,\DSP_PREADD_DATA.A2A1<24> ,\DSP_PREADD_DATA.A2A1<23> ,\DSP_PREADD_DATA.A2A1<22> ,\DSP_PREADD_DATA.A2A1<21> ,\DSP_PREADD_DATA.A2A1<20> ,\DSP_PREADD_DATA.A2A1<19> ,\DSP_PREADD_DATA.A2A1<18> ,\DSP_PREADD_DATA.A2A1<17> ,\DSP_PREADD_DATA.A2A1<16> ,\DSP_PREADD_DATA.A2A1<15> ,\DSP_PREADD_DATA.A2A1<14> ,\DSP_PREADD_DATA.A2A1<13> ,\DSP_PREADD_DATA.A2A1<12> ,\DSP_PREADD_DATA.A2A1<11> ,\DSP_PREADD_DATA.A2A1<10> ,\DSP_PREADD_DATA.A2A1<9> ,\DSP_PREADD_DATA.A2A1<8> ,\DSP_PREADD_DATA.A2A1<7> ,\DSP_PREADD_DATA.A2A1<6> ,\DSP_PREADD_DATA.A2A1<5> ,\DSP_PREADD_DATA.A2A1<4> ,\DSP_PREADD_DATA.A2A1<3> ,\DSP_PREADD_DATA.A2A1<2> ,\DSP_PREADD_DATA.A2A1<1> ,\DSP_PREADD_DATA.A2A1<0> }),
        .AD_DATA({\DSP_PREADD_DATA.AD_DATA<26> ,\DSP_PREADD_DATA.AD_DATA<25> ,\DSP_PREADD_DATA.AD_DATA<24> ,\DSP_PREADD_DATA.AD_DATA<23> ,\DSP_PREADD_DATA.AD_DATA<22> ,\DSP_PREADD_DATA.AD_DATA<21> ,\DSP_PREADD_DATA.AD_DATA<20> ,\DSP_PREADD_DATA.AD_DATA<19> ,\DSP_PREADD_DATA.AD_DATA<18> ,\DSP_PREADD_DATA.AD_DATA<17> ,\DSP_PREADD_DATA.AD_DATA<16> ,\DSP_PREADD_DATA.AD_DATA<15> ,\DSP_PREADD_DATA.AD_DATA<14> ,\DSP_PREADD_DATA.AD_DATA<13> ,\DSP_PREADD_DATA.AD_DATA<12> ,\DSP_PREADD_DATA.AD_DATA<11> ,\DSP_PREADD_DATA.AD_DATA<10> ,\DSP_PREADD_DATA.AD_DATA<9> ,\DSP_PREADD_DATA.AD_DATA<8> ,\DSP_PREADD_DATA.AD_DATA<7> ,\DSP_PREADD_DATA.AD_DATA<6> ,\DSP_PREADD_DATA.AD_DATA<5> ,\DSP_PREADD_DATA.AD_DATA<4> ,\DSP_PREADD_DATA.AD_DATA<3> ,\DSP_PREADD_DATA.AD_DATA<2> ,\DSP_PREADD_DATA.AD_DATA<1> ,\DSP_PREADD_DATA.AD_DATA<0> }),
        .AMULT26(\DSP_MULTIPLIER.AMULT26 ),
        .B2B1({\DSP_PREADD_DATA.B2B1<17> ,\DSP_PREADD_DATA.B2B1<16> ,\DSP_PREADD_DATA.B2B1<15> ,\DSP_PREADD_DATA.B2B1<14> ,\DSP_PREADD_DATA.B2B1<13> ,\DSP_PREADD_DATA.B2B1<12> ,\DSP_PREADD_DATA.B2B1<11> ,\DSP_PREADD_DATA.B2B1<10> ,\DSP_PREADD_DATA.B2B1<9> ,\DSP_PREADD_DATA.B2B1<8> ,\DSP_PREADD_DATA.B2B1<7> ,\DSP_PREADD_DATA.B2B1<6> ,\DSP_PREADD_DATA.B2B1<5> ,\DSP_PREADD_DATA.B2B1<4> ,\DSP_PREADD_DATA.B2B1<3> ,\DSP_PREADD_DATA.B2B1<2> ,\DSP_PREADD_DATA.B2B1<1> ,\DSP_PREADD_DATA.B2B1<0> }),
        .BMULT17(\DSP_MULTIPLIER.BMULT17 ),
        .U({\DSP_MULTIPLIER.U<44> ,\DSP_MULTIPLIER.U<43> ,\DSP_MULTIPLIER.U<42> ,\DSP_MULTIPLIER.U<41> ,\DSP_MULTIPLIER.U<40> ,\DSP_MULTIPLIER.U<39> ,\DSP_MULTIPLIER.U<38> ,\DSP_MULTIPLIER.U<37> ,\DSP_MULTIPLIER.U<36> ,\DSP_MULTIPLIER.U<35> ,\DSP_MULTIPLIER.U<34> ,\DSP_MULTIPLIER.U<33> ,\DSP_MULTIPLIER.U<32> ,\DSP_MULTIPLIER.U<31> ,\DSP_MULTIPLIER.U<30> ,\DSP_MULTIPLIER.U<29> ,\DSP_MULTIPLIER.U<28> ,\DSP_MULTIPLIER.U<27> ,\DSP_MULTIPLIER.U<26> ,\DSP_MULTIPLIER.U<25> ,\DSP_MULTIPLIER.U<24> ,\DSP_MULTIPLIER.U<23> ,\DSP_MULTIPLIER.U<22> ,\DSP_MULTIPLIER.U<21> ,\DSP_MULTIPLIER.U<20> ,\DSP_MULTIPLIER.U<19> ,\DSP_MULTIPLIER.U<18> ,\DSP_MULTIPLIER.U<17> ,\DSP_MULTIPLIER.U<16> ,\DSP_MULTIPLIER.U<15> ,\DSP_MULTIPLIER.U<14> ,\DSP_MULTIPLIER.U<13> ,\DSP_MULTIPLIER.U<12> ,\DSP_MULTIPLIER.U<11> ,\DSP_MULTIPLIER.U<10> ,\DSP_MULTIPLIER.U<9> ,\DSP_MULTIPLIER.U<8> ,\DSP_MULTIPLIER.U<7> ,\DSP_MULTIPLIER.U<6> ,\DSP_MULTIPLIER.U<5> ,\DSP_MULTIPLIER.U<4> ,\DSP_MULTIPLIER.U<3> ,\DSP_MULTIPLIER.U<2> ,\DSP_MULTIPLIER.U<1> ,\DSP_MULTIPLIER.U<0> }),
        .V({\DSP_MULTIPLIER.V<44> ,\DSP_MULTIPLIER.V<43> ,\DSP_MULTIPLIER.V<42> ,\DSP_MULTIPLIER.V<41> ,\DSP_MULTIPLIER.V<40> ,\DSP_MULTIPLIER.V<39> ,\DSP_MULTIPLIER.V<38> ,\DSP_MULTIPLIER.V<37> ,\DSP_MULTIPLIER.V<36> ,\DSP_MULTIPLIER.V<35> ,\DSP_MULTIPLIER.V<34> ,\DSP_MULTIPLIER.V<33> ,\DSP_MULTIPLIER.V<32> ,\DSP_MULTIPLIER.V<31> ,\DSP_MULTIPLIER.V<30> ,\DSP_MULTIPLIER.V<29> ,\DSP_MULTIPLIER.V<28> ,\DSP_MULTIPLIER.V<27> ,\DSP_MULTIPLIER.V<26> ,\DSP_MULTIPLIER.V<25> ,\DSP_MULTIPLIER.V<24> ,\DSP_MULTIPLIER.V<23> ,\DSP_MULTIPLIER.V<22> ,\DSP_MULTIPLIER.V<21> ,\DSP_MULTIPLIER.V<20> ,\DSP_MULTIPLIER.V<19> ,\DSP_MULTIPLIER.V<18> ,\DSP_MULTIPLIER.V<17> ,\DSP_MULTIPLIER.V<16> ,\DSP_MULTIPLIER.V<15> ,\DSP_MULTIPLIER.V<14> ,\DSP_MULTIPLIER.V<13> ,\DSP_MULTIPLIER.V<12> ,\DSP_MULTIPLIER.V<11> ,\DSP_MULTIPLIER.V<10> ,\DSP_MULTIPLIER.V<9> ,\DSP_MULTIPLIER.V<8> ,\DSP_MULTIPLIER.V<7> ,\DSP_MULTIPLIER.V<6> ,\DSP_MULTIPLIER.V<5> ,\DSP_MULTIPLIER.V<4> ,\DSP_MULTIPLIER.V<3> ,\DSP_MULTIPLIER.V<2> ,\DSP_MULTIPLIER.V<1> ,\DSP_MULTIPLIER.V<0> }));
  DSP_M_DATA #(
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .MREG(0)) 
    DSP_M_DATA_INST
       (.CEM(CEM),
        .CLK(CLK),
        .RSTM(RSTM),
        .U({\DSP_MULTIPLIER.U<44> ,\DSP_MULTIPLIER.U<43> ,\DSP_MULTIPLIER.U<42> ,\DSP_MULTIPLIER.U<41> ,\DSP_MULTIPLIER.U<40> ,\DSP_MULTIPLIER.U<39> ,\DSP_MULTIPLIER.U<38> ,\DSP_MULTIPLIER.U<37> ,\DSP_MULTIPLIER.U<36> ,\DSP_MULTIPLIER.U<35> ,\DSP_MULTIPLIER.U<34> ,\DSP_MULTIPLIER.U<33> ,\DSP_MULTIPLIER.U<32> ,\DSP_MULTIPLIER.U<31> ,\DSP_MULTIPLIER.U<30> ,\DSP_MULTIPLIER.U<29> ,\DSP_MULTIPLIER.U<28> ,\DSP_MULTIPLIER.U<27> ,\DSP_MULTIPLIER.U<26> ,\DSP_MULTIPLIER.U<25> ,\DSP_MULTIPLIER.U<24> ,\DSP_MULTIPLIER.U<23> ,\DSP_MULTIPLIER.U<22> ,\DSP_MULTIPLIER.U<21> ,\DSP_MULTIPLIER.U<20> ,\DSP_MULTIPLIER.U<19> ,\DSP_MULTIPLIER.U<18> ,\DSP_MULTIPLIER.U<17> ,\DSP_MULTIPLIER.U<16> ,\DSP_MULTIPLIER.U<15> ,\DSP_MULTIPLIER.U<14> ,\DSP_MULTIPLIER.U<13> ,\DSP_MULTIPLIER.U<12> ,\DSP_MULTIPLIER.U<11> ,\DSP_MULTIPLIER.U<10> ,\DSP_MULTIPLIER.U<9> ,\DSP_MULTIPLIER.U<8> ,\DSP_MULTIPLIER.U<7> ,\DSP_MULTIPLIER.U<6> ,\DSP_MULTIPLIER.U<5> ,\DSP_MULTIPLIER.U<4> ,\DSP_MULTIPLIER.U<3> ,\DSP_MULTIPLIER.U<2> ,\DSP_MULTIPLIER.U<1> ,\DSP_MULTIPLIER.U<0> }),
        .U_DATA({\DSP_M_DATA.U_DATA<44> ,\DSP_M_DATA.U_DATA<43> ,\DSP_M_DATA.U_DATA<42> ,\DSP_M_DATA.U_DATA<41> ,\DSP_M_DATA.U_DATA<40> ,\DSP_M_DATA.U_DATA<39> ,\DSP_M_DATA.U_DATA<38> ,\DSP_M_DATA.U_DATA<37> ,\DSP_M_DATA.U_DATA<36> ,\DSP_M_DATA.U_DATA<35> ,\DSP_M_DATA.U_DATA<34> ,\DSP_M_DATA.U_DATA<33> ,\DSP_M_DATA.U_DATA<32> ,\DSP_M_DATA.U_DATA<31> ,\DSP_M_DATA.U_DATA<30> ,\DSP_M_DATA.U_DATA<29> ,\DSP_M_DATA.U_DATA<28> ,\DSP_M_DATA.U_DATA<27> ,\DSP_M_DATA.U_DATA<26> ,\DSP_M_DATA.U_DATA<25> ,\DSP_M_DATA.U_DATA<24> ,\DSP_M_DATA.U_DATA<23> ,\DSP_M_DATA.U_DATA<22> ,\DSP_M_DATA.U_DATA<21> ,\DSP_M_DATA.U_DATA<20> ,\DSP_M_DATA.U_DATA<19> ,\DSP_M_DATA.U_DATA<18> ,\DSP_M_DATA.U_DATA<17> ,\DSP_M_DATA.U_DATA<16> ,\DSP_M_DATA.U_DATA<15> ,\DSP_M_DATA.U_DATA<14> ,\DSP_M_DATA.U_DATA<13> ,\DSP_M_DATA.U_DATA<12> ,\DSP_M_DATA.U_DATA<11> ,\DSP_M_DATA.U_DATA<10> ,\DSP_M_DATA.U_DATA<9> ,\DSP_M_DATA.U_DATA<8> ,\DSP_M_DATA.U_DATA<7> ,\DSP_M_DATA.U_DATA<6> ,\DSP_M_DATA.U_DATA<5> ,\DSP_M_DATA.U_DATA<4> ,\DSP_M_DATA.U_DATA<3> ,\DSP_M_DATA.U_DATA<2> ,\DSP_M_DATA.U_DATA<1> ,\DSP_M_DATA.U_DATA<0> }),
        .V({\DSP_MULTIPLIER.V<44> ,\DSP_MULTIPLIER.V<43> ,\DSP_MULTIPLIER.V<42> ,\DSP_MULTIPLIER.V<41> ,\DSP_MULTIPLIER.V<40> ,\DSP_MULTIPLIER.V<39> ,\DSP_MULTIPLIER.V<38> ,\DSP_MULTIPLIER.V<37> ,\DSP_MULTIPLIER.V<36> ,\DSP_MULTIPLIER.V<35> ,\DSP_MULTIPLIER.V<34> ,\DSP_MULTIPLIER.V<33> ,\DSP_MULTIPLIER.V<32> ,\DSP_MULTIPLIER.V<31> ,\DSP_MULTIPLIER.V<30> ,\DSP_MULTIPLIER.V<29> ,\DSP_MULTIPLIER.V<28> ,\DSP_MULTIPLIER.V<27> ,\DSP_MULTIPLIER.V<26> ,\DSP_MULTIPLIER.V<25> ,\DSP_MULTIPLIER.V<24> ,\DSP_MULTIPLIER.V<23> ,\DSP_MULTIPLIER.V<22> ,\DSP_MULTIPLIER.V<21> ,\DSP_MULTIPLIER.V<20> ,\DSP_MULTIPLIER.V<19> ,\DSP_MULTIPLIER.V<18> ,\DSP_MULTIPLIER.V<17> ,\DSP_MULTIPLIER.V<16> ,\DSP_MULTIPLIER.V<15> ,\DSP_MULTIPLIER.V<14> ,\DSP_MULTIPLIER.V<13> ,\DSP_MULTIPLIER.V<12> ,\DSP_MULTIPLIER.V<11> ,\DSP_MULTIPLIER.V<10> ,\DSP_MULTIPLIER.V<9> ,\DSP_MULTIPLIER.V<8> ,\DSP_MULTIPLIER.V<7> ,\DSP_MULTIPLIER.V<6> ,\DSP_MULTIPLIER.V<5> ,\DSP_MULTIPLIER.V<4> ,\DSP_MULTIPLIER.V<3> ,\DSP_MULTIPLIER.V<2> ,\DSP_MULTIPLIER.V<1> ,\DSP_MULTIPLIER.V<0> }),
        .V_DATA({\DSP_M_DATA.V_DATA<44> ,\DSP_M_DATA.V_DATA<43> ,\DSP_M_DATA.V_DATA<42> ,\DSP_M_DATA.V_DATA<41> ,\DSP_M_DATA.V_DATA<40> ,\DSP_M_DATA.V_DATA<39> ,\DSP_M_DATA.V_DATA<38> ,\DSP_M_DATA.V_DATA<37> ,\DSP_M_DATA.V_DATA<36> ,\DSP_M_DATA.V_DATA<35> ,\DSP_M_DATA.V_DATA<34> ,\DSP_M_DATA.V_DATA<33> ,\DSP_M_DATA.V_DATA<32> ,\DSP_M_DATA.V_DATA<31> ,\DSP_M_DATA.V_DATA<30> ,\DSP_M_DATA.V_DATA<29> ,\DSP_M_DATA.V_DATA<28> ,\DSP_M_DATA.V_DATA<27> ,\DSP_M_DATA.V_DATA<26> ,\DSP_M_DATA.V_DATA<25> ,\DSP_M_DATA.V_DATA<24> ,\DSP_M_DATA.V_DATA<23> ,\DSP_M_DATA.V_DATA<22> ,\DSP_M_DATA.V_DATA<21> ,\DSP_M_DATA.V_DATA<20> ,\DSP_M_DATA.V_DATA<19> ,\DSP_M_DATA.V_DATA<18> ,\DSP_M_DATA.V_DATA<17> ,\DSP_M_DATA.V_DATA<16> ,\DSP_M_DATA.V_DATA<15> ,\DSP_M_DATA.V_DATA<14> ,\DSP_M_DATA.V_DATA<13> ,\DSP_M_DATA.V_DATA<12> ,\DSP_M_DATA.V_DATA<11> ,\DSP_M_DATA.V_DATA<10> ,\DSP_M_DATA.V_DATA<9> ,\DSP_M_DATA.V_DATA<8> ,\DSP_M_DATA.V_DATA<7> ,\DSP_M_DATA.V_DATA<6> ,\DSP_M_DATA.V_DATA<5> ,\DSP_M_DATA.V_DATA<4> ,\DSP_M_DATA.V_DATA<3> ,\DSP_M_DATA.V_DATA<2> ,\DSP_M_DATA.V_DATA<1> ,\DSP_M_DATA.V_DATA<0> }));
  DSP_OUTPUT #(
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .IS_CLK_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h3FFFFFFFFFFF),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_PATTERN_DETECT("NO_PATDET")) 
    DSP_OUTPUT_INST
       (.ALUMODE10(\DSP_ALU.ALUMODE10 ),
        .ALU_OUT({\DSP_ALU.ALU_OUT<47> ,\DSP_ALU.ALU_OUT<46> ,\DSP_ALU.ALU_OUT<45> ,\DSP_ALU.ALU_OUT<44> ,\DSP_ALU.ALU_OUT<43> ,\DSP_ALU.ALU_OUT<42> ,\DSP_ALU.ALU_OUT<41> ,\DSP_ALU.ALU_OUT<40> ,\DSP_ALU.ALU_OUT<39> ,\DSP_ALU.ALU_OUT<38> ,\DSP_ALU.ALU_OUT<37> ,\DSP_ALU.ALU_OUT<36> ,\DSP_ALU.ALU_OUT<35> ,\DSP_ALU.ALU_OUT<34> ,\DSP_ALU.ALU_OUT<33> ,\DSP_ALU.ALU_OUT<32> ,\DSP_ALU.ALU_OUT<31> ,\DSP_ALU.ALU_OUT<30> ,\DSP_ALU.ALU_OUT<29> ,\DSP_ALU.ALU_OUT<28> ,\DSP_ALU.ALU_OUT<27> ,\DSP_ALU.ALU_OUT<26> ,\DSP_ALU.ALU_OUT<25> ,\DSP_ALU.ALU_OUT<24> ,\DSP_ALU.ALU_OUT<23> ,\DSP_ALU.ALU_OUT<22> ,\DSP_ALU.ALU_OUT<21> ,\DSP_ALU.ALU_OUT<20> ,\DSP_ALU.ALU_OUT<19> ,\DSP_ALU.ALU_OUT<18> ,\DSP_ALU.ALU_OUT<17> ,\DSP_ALU.ALU_OUT<16> ,\DSP_ALU.ALU_OUT<15> ,\DSP_ALU.ALU_OUT<14> ,\DSP_ALU.ALU_OUT<13> ,\DSP_ALU.ALU_OUT<12> ,\DSP_ALU.ALU_OUT<11> ,\DSP_ALU.ALU_OUT<10> ,\DSP_ALU.ALU_OUT<9> ,\DSP_ALU.ALU_OUT<8> ,\DSP_ALU.ALU_OUT<7> ,\DSP_ALU.ALU_OUT<6> ,\DSP_ALU.ALU_OUT<5> ,\DSP_ALU.ALU_OUT<4> ,\DSP_ALU.ALU_OUT<3> ,\DSP_ALU.ALU_OUT<2> ,\DSP_ALU.ALU_OUT<1> ,\DSP_ALU.ALU_OUT<0> }),
        .CARRYCASCOUT(CARRYCASCOUT),
        .CARRYOUT({\CARRYOUT[3] ,\CARRYOUT[2] ,\CARRYOUT[1] ,\CARRYOUT[0] }),
        .CCOUT_FB(\DSP_OUTPUT.CCOUT_FB ),
        .CEP(CEP),
        .CLK(CLK),
        .COUT({\DSP_ALU.COUT<3> ,\DSP_ALU.COUT<2> ,\DSP_ALU.COUT<1> ,\DSP_ALU.COUT<0> }),
        .C_DATA({\DSP_C_DATA.C_DATA<47> ,\DSP_C_DATA.C_DATA<46> ,\DSP_C_DATA.C_DATA<45> ,\DSP_C_DATA.C_DATA<44> ,\DSP_C_DATA.C_DATA<43> ,\DSP_C_DATA.C_DATA<42> ,\DSP_C_DATA.C_DATA<41> ,\DSP_C_DATA.C_DATA<40> ,\DSP_C_DATA.C_DATA<39> ,\DSP_C_DATA.C_DATA<38> ,\DSP_C_DATA.C_DATA<37> ,\DSP_C_DATA.C_DATA<36> ,\DSP_C_DATA.C_DATA<35> ,\DSP_C_DATA.C_DATA<34> ,\DSP_C_DATA.C_DATA<33> ,\DSP_C_DATA.C_DATA<32> ,\DSP_C_DATA.C_DATA<31> ,\DSP_C_DATA.C_DATA<30> ,\DSP_C_DATA.C_DATA<29> ,\DSP_C_DATA.C_DATA<28> ,\DSP_C_DATA.C_DATA<27> ,\DSP_C_DATA.C_DATA<26> ,\DSP_C_DATA.C_DATA<25> ,\DSP_C_DATA.C_DATA<24> ,\DSP_C_DATA.C_DATA<23> ,\DSP_C_DATA.C_DATA<22> ,\DSP_C_DATA.C_DATA<21> ,\DSP_C_DATA.C_DATA<20> ,\DSP_C_DATA.C_DATA<19> ,\DSP_C_DATA.C_DATA<18> ,\DSP_C_DATA.C_DATA<17> ,\DSP_C_DATA.C_DATA<16> ,\DSP_C_DATA.C_DATA<15> ,\DSP_C_DATA.C_DATA<14> ,\DSP_C_DATA.C_DATA<13> ,\DSP_C_DATA.C_DATA<12> ,\DSP_C_DATA.C_DATA<11> ,\DSP_C_DATA.C_DATA<10> ,\DSP_C_DATA.C_DATA<9> ,\DSP_C_DATA.C_DATA<8> ,\DSP_C_DATA.C_DATA<7> ,\DSP_C_DATA.C_DATA<6> ,\DSP_C_DATA.C_DATA<5> ,\DSP_C_DATA.C_DATA<4> ,\DSP_C_DATA.C_DATA<3> ,\DSP_C_DATA.C_DATA<2> ,\DSP_C_DATA.C_DATA<1> ,\DSP_C_DATA.C_DATA<0> }),
        .MULTSIGNOUT(MULTSIGNOUT),
        .MULTSIGN_ALU(\DSP_ALU.MULTSIGN_ALU ),
        .OVERFLOW(OVERFLOW),
        .P({\P[47] ,\P[46] ,\P[45] ,\P[44] ,\P[43] ,\P[42] ,\P[41] ,\P[40] ,\P[39] ,\P[38] ,\P[37] ,\P[36] ,\P[35] ,\P[34] ,\P[33] ,\P[32] ,\P[31] ,\P[30] ,\P[29] ,\P[28] ,\P[27] ,\P[26] ,\P[25] ,\P[24] ,\P[23] ,\P[22] ,\P[21] ,\P[20] ,\P[19] ,\P[18] ,\P[17] ,\P[16] ,\P[15] ,\P[14] ,\P[13] ,\P[12] ,\P[11] ,\P[10] ,\P[9] ,\P[8] ,\P[7] ,\P[6] ,\P[5] ,\P[4] ,\P[3] ,\P[2] ,\P[1] ,\P[0] }),
        .PATTERN_B_DETECT(PATTERNBDETECT),
        .PATTERN_DETECT(PATTERNDETECT),
        .PCOUT({\PCOUT[47] ,\PCOUT[46] ,\PCOUT[45] ,\PCOUT[44] ,\PCOUT[43] ,\PCOUT[42] ,\PCOUT[41] ,\PCOUT[40] ,\PCOUT[39] ,\PCOUT[38] ,\PCOUT[37] ,\PCOUT[36] ,\PCOUT[35] ,\PCOUT[34] ,\PCOUT[33] ,\PCOUT[32] ,\PCOUT[31] ,\PCOUT[30] ,\PCOUT[29] ,\PCOUT[28] ,\PCOUT[27] ,\PCOUT[26] ,\PCOUT[25] ,\PCOUT[24] ,\PCOUT[23] ,\PCOUT[22] ,\PCOUT[21] ,\PCOUT[20] ,\PCOUT[19] ,\PCOUT[18] ,\PCOUT[17] ,\PCOUT[16] ,\PCOUT[15] ,\PCOUT[14] ,\PCOUT[13] ,\PCOUT[12] ,\PCOUT[11] ,\PCOUT[10] ,\PCOUT[9] ,\PCOUT[8] ,\PCOUT[7] ,\PCOUT[6] ,\PCOUT[5] ,\PCOUT[4] ,\PCOUT[3] ,\PCOUT[2] ,\PCOUT[1] ,\PCOUT[0] }),
        .P_FDBK({\DSP_OUTPUT.P_FDBK<47> ,\DSP_OUTPUT.P_FDBK<46> ,\DSP_OUTPUT.P_FDBK<45> ,\DSP_OUTPUT.P_FDBK<44> ,\DSP_OUTPUT.P_FDBK<43> ,\DSP_OUTPUT.P_FDBK<42> ,\DSP_OUTPUT.P_FDBK<41> ,\DSP_OUTPUT.P_FDBK<40> ,\DSP_OUTPUT.P_FDBK<39> ,\DSP_OUTPUT.P_FDBK<38> ,\DSP_OUTPUT.P_FDBK<37> ,\DSP_OUTPUT.P_FDBK<36> ,\DSP_OUTPUT.P_FDBK<35> ,\DSP_OUTPUT.P_FDBK<34> ,\DSP_OUTPUT.P_FDBK<33> ,\DSP_OUTPUT.P_FDBK<32> ,\DSP_OUTPUT.P_FDBK<31> ,\DSP_OUTPUT.P_FDBK<30> ,\DSP_OUTPUT.P_FDBK<29> ,\DSP_OUTPUT.P_FDBK<28> ,\DSP_OUTPUT.P_FDBK<27> ,\DSP_OUTPUT.P_FDBK<26> ,\DSP_OUTPUT.P_FDBK<25> ,\DSP_OUTPUT.P_FDBK<24> ,\DSP_OUTPUT.P_FDBK<23> ,\DSP_OUTPUT.P_FDBK<22> ,\DSP_OUTPUT.P_FDBK<21> ,\DSP_OUTPUT.P_FDBK<20> ,\DSP_OUTPUT.P_FDBK<19> ,\DSP_OUTPUT.P_FDBK<18> ,\DSP_OUTPUT.P_FDBK<17> ,\DSP_OUTPUT.P_FDBK<16> ,\DSP_OUTPUT.P_FDBK<15> ,\DSP_OUTPUT.P_FDBK<14> ,\DSP_OUTPUT.P_FDBK<13> ,\DSP_OUTPUT.P_FDBK<12> ,\DSP_OUTPUT.P_FDBK<11> ,\DSP_OUTPUT.P_FDBK<10> ,\DSP_OUTPUT.P_FDBK<9> ,\DSP_OUTPUT.P_FDBK<8> ,\DSP_OUTPUT.P_FDBK<7> ,\DSP_OUTPUT.P_FDBK<6> ,\DSP_OUTPUT.P_FDBK<5> ,\DSP_OUTPUT.P_FDBK<4> ,\DSP_OUTPUT.P_FDBK<3> ,\DSP_OUTPUT.P_FDBK<2> ,\DSP_OUTPUT.P_FDBK<1> ,\DSP_OUTPUT.P_FDBK<0> }),
        .P_FDBK_47(\DSP_OUTPUT.P_FDBK_47 ),
        .RSTP(RSTP),
        .UNDERFLOW(UNDERFLOW),
        .XOROUT({\XOROUT[7] ,\XOROUT[6] ,\XOROUT[5] ,\XOROUT[4] ,\XOROUT[3] ,\XOROUT[2] ,\XOROUT[1] ,\XOROUT[0] }),
        .XOR_MX({\DSP_ALU.XOR_MX<7> ,\DSP_ALU.XOR_MX<6> ,\DSP_ALU.XOR_MX<5> ,\DSP_ALU.XOR_MX<4> ,\DSP_ALU.XOR_MX<3> ,\DSP_ALU.XOR_MX<2> ,\DSP_ALU.XOR_MX<1> ,\DSP_ALU.XOR_MX<0> }));
  DSP_PREADD_DATA #(
    .ADREG(1),
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .DREG(1),
    .INMODEREG(0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .PREADDINSEL("A"),
    .USE_MULT("MULTIPLY")) 
    DSP_PREADD_DATA_INST
       (.A1_DATA({\DSP_A_B_DATA.A1_DATA<26> ,\DSP_A_B_DATA.A1_DATA<25> ,\DSP_A_B_DATA.A1_DATA<24> ,\DSP_A_B_DATA.A1_DATA<23> ,\DSP_A_B_DATA.A1_DATA<22> ,\DSP_A_B_DATA.A1_DATA<21> ,\DSP_A_B_DATA.A1_DATA<20> ,\DSP_A_B_DATA.A1_DATA<19> ,\DSP_A_B_DATA.A1_DATA<18> ,\DSP_A_B_DATA.A1_DATA<17> ,\DSP_A_B_DATA.A1_DATA<16> ,\DSP_A_B_DATA.A1_DATA<15> ,\DSP_A_B_DATA.A1_DATA<14> ,\DSP_A_B_DATA.A1_DATA<13> ,\DSP_A_B_DATA.A1_DATA<12> ,\DSP_A_B_DATA.A1_DATA<11> ,\DSP_A_B_DATA.A1_DATA<10> ,\DSP_A_B_DATA.A1_DATA<9> ,\DSP_A_B_DATA.A1_DATA<8> ,\DSP_A_B_DATA.A1_DATA<7> ,\DSP_A_B_DATA.A1_DATA<6> ,\DSP_A_B_DATA.A1_DATA<5> ,\DSP_A_B_DATA.A1_DATA<4> ,\DSP_A_B_DATA.A1_DATA<3> ,\DSP_A_B_DATA.A1_DATA<2> ,\DSP_A_B_DATA.A1_DATA<1> ,\DSP_A_B_DATA.A1_DATA<0> }),
        .A2A1({\DSP_PREADD_DATA.A2A1<26> ,\DSP_PREADD_DATA.A2A1<25> ,\DSP_PREADD_DATA.A2A1<24> ,\DSP_PREADD_DATA.A2A1<23> ,\DSP_PREADD_DATA.A2A1<22> ,\DSP_PREADD_DATA.A2A1<21> ,\DSP_PREADD_DATA.A2A1<20> ,\DSP_PREADD_DATA.A2A1<19> ,\DSP_PREADD_DATA.A2A1<18> ,\DSP_PREADD_DATA.A2A1<17> ,\DSP_PREADD_DATA.A2A1<16> ,\DSP_PREADD_DATA.A2A1<15> ,\DSP_PREADD_DATA.A2A1<14> ,\DSP_PREADD_DATA.A2A1<13> ,\DSP_PREADD_DATA.A2A1<12> ,\DSP_PREADD_DATA.A2A1<11> ,\DSP_PREADD_DATA.A2A1<10> ,\DSP_PREADD_DATA.A2A1<9> ,\DSP_PREADD_DATA.A2A1<8> ,\DSP_PREADD_DATA.A2A1<7> ,\DSP_PREADD_DATA.A2A1<6> ,\DSP_PREADD_DATA.A2A1<5> ,\DSP_PREADD_DATA.A2A1<4> ,\DSP_PREADD_DATA.A2A1<3> ,\DSP_PREADD_DATA.A2A1<2> ,\DSP_PREADD_DATA.A2A1<1> ,\DSP_PREADD_DATA.A2A1<0> }),
        .A2_DATA({\DSP_A_B_DATA.A2_DATA<26> ,\DSP_A_B_DATA.A2_DATA<25> ,\DSP_A_B_DATA.A2_DATA<24> ,\DSP_A_B_DATA.A2_DATA<23> ,\DSP_A_B_DATA.A2_DATA<22> ,\DSP_A_B_DATA.A2_DATA<21> ,\DSP_A_B_DATA.A2_DATA<20> ,\DSP_A_B_DATA.A2_DATA<19> ,\DSP_A_B_DATA.A2_DATA<18> ,\DSP_A_B_DATA.A2_DATA<17> ,\DSP_A_B_DATA.A2_DATA<16> ,\DSP_A_B_DATA.A2_DATA<15> ,\DSP_A_B_DATA.A2_DATA<14> ,\DSP_A_B_DATA.A2_DATA<13> ,\DSP_A_B_DATA.A2_DATA<12> ,\DSP_A_B_DATA.A2_DATA<11> ,\DSP_A_B_DATA.A2_DATA<10> ,\DSP_A_B_DATA.A2_DATA<9> ,\DSP_A_B_DATA.A2_DATA<8> ,\DSP_A_B_DATA.A2_DATA<7> ,\DSP_A_B_DATA.A2_DATA<6> ,\DSP_A_B_DATA.A2_DATA<5> ,\DSP_A_B_DATA.A2_DATA<4> ,\DSP_A_B_DATA.A2_DATA<3> ,\DSP_A_B_DATA.A2_DATA<2> ,\DSP_A_B_DATA.A2_DATA<1> ,\DSP_A_B_DATA.A2_DATA<0> }),
        .AD({\DSP_PREADD.AD<26> ,\DSP_PREADD.AD<25> ,\DSP_PREADD.AD<24> ,\DSP_PREADD.AD<23> ,\DSP_PREADD.AD<22> ,\DSP_PREADD.AD<21> ,\DSP_PREADD.AD<20> ,\DSP_PREADD.AD<19> ,\DSP_PREADD.AD<18> ,\DSP_PREADD.AD<17> ,\DSP_PREADD.AD<16> ,\DSP_PREADD.AD<15> ,\DSP_PREADD.AD<14> ,\DSP_PREADD.AD<13> ,\DSP_PREADD.AD<12> ,\DSP_PREADD.AD<11> ,\DSP_PREADD.AD<10> ,\DSP_PREADD.AD<9> ,\DSP_PREADD.AD<8> ,\DSP_PREADD.AD<7> ,\DSP_PREADD.AD<6> ,\DSP_PREADD.AD<5> ,\DSP_PREADD.AD<4> ,\DSP_PREADD.AD<3> ,\DSP_PREADD.AD<2> ,\DSP_PREADD.AD<1> ,\DSP_PREADD.AD<0> }),
        .ADDSUB(\DSP_PREADD_DATA.ADDSUB ),
        .AD_DATA({\DSP_PREADD_DATA.AD_DATA<26> ,\DSP_PREADD_DATA.AD_DATA<25> ,\DSP_PREADD_DATA.AD_DATA<24> ,\DSP_PREADD_DATA.AD_DATA<23> ,\DSP_PREADD_DATA.AD_DATA<22> ,\DSP_PREADD_DATA.AD_DATA<21> ,\DSP_PREADD_DATA.AD_DATA<20> ,\DSP_PREADD_DATA.AD_DATA<19> ,\DSP_PREADD_DATA.AD_DATA<18> ,\DSP_PREADD_DATA.AD_DATA<17> ,\DSP_PREADD_DATA.AD_DATA<16> ,\DSP_PREADD_DATA.AD_DATA<15> ,\DSP_PREADD_DATA.AD_DATA<14> ,\DSP_PREADD_DATA.AD_DATA<13> ,\DSP_PREADD_DATA.AD_DATA<12> ,\DSP_PREADD_DATA.AD_DATA<11> ,\DSP_PREADD_DATA.AD_DATA<10> ,\DSP_PREADD_DATA.AD_DATA<9> ,\DSP_PREADD_DATA.AD_DATA<8> ,\DSP_PREADD_DATA.AD_DATA<7> ,\DSP_PREADD_DATA.AD_DATA<6> ,\DSP_PREADD_DATA.AD_DATA<5> ,\DSP_PREADD_DATA.AD_DATA<4> ,\DSP_PREADD_DATA.AD_DATA<3> ,\DSP_PREADD_DATA.AD_DATA<2> ,\DSP_PREADD_DATA.AD_DATA<1> ,\DSP_PREADD_DATA.AD_DATA<0> }),
        .B1_DATA({\DSP_A_B_DATA.B1_DATA<17> ,\DSP_A_B_DATA.B1_DATA<16> ,\DSP_A_B_DATA.B1_DATA<15> ,\DSP_A_B_DATA.B1_DATA<14> ,\DSP_A_B_DATA.B1_DATA<13> ,\DSP_A_B_DATA.B1_DATA<12> ,\DSP_A_B_DATA.B1_DATA<11> ,\DSP_A_B_DATA.B1_DATA<10> ,\DSP_A_B_DATA.B1_DATA<9> ,\DSP_A_B_DATA.B1_DATA<8> ,\DSP_A_B_DATA.B1_DATA<7> ,\DSP_A_B_DATA.B1_DATA<6> ,\DSP_A_B_DATA.B1_DATA<5> ,\DSP_A_B_DATA.B1_DATA<4> ,\DSP_A_B_DATA.B1_DATA<3> ,\DSP_A_B_DATA.B1_DATA<2> ,\DSP_A_B_DATA.B1_DATA<1> ,\DSP_A_B_DATA.B1_DATA<0> }),
        .B2B1({\DSP_PREADD_DATA.B2B1<17> ,\DSP_PREADD_DATA.B2B1<16> ,\DSP_PREADD_DATA.B2B1<15> ,\DSP_PREADD_DATA.B2B1<14> ,\DSP_PREADD_DATA.B2B1<13> ,\DSP_PREADD_DATA.B2B1<12> ,\DSP_PREADD_DATA.B2B1<11> ,\DSP_PREADD_DATA.B2B1<10> ,\DSP_PREADD_DATA.B2B1<9> ,\DSP_PREADD_DATA.B2B1<8> ,\DSP_PREADD_DATA.B2B1<7> ,\DSP_PREADD_DATA.B2B1<6> ,\DSP_PREADD_DATA.B2B1<5> ,\DSP_PREADD_DATA.B2B1<4> ,\DSP_PREADD_DATA.B2B1<3> ,\DSP_PREADD_DATA.B2B1<2> ,\DSP_PREADD_DATA.B2B1<1> ,\DSP_PREADD_DATA.B2B1<0> }),
        .B2_DATA({\DSP_A_B_DATA.B2_DATA<17> ,\DSP_A_B_DATA.B2_DATA<16> ,\DSP_A_B_DATA.B2_DATA<15> ,\DSP_A_B_DATA.B2_DATA<14> ,\DSP_A_B_DATA.B2_DATA<13> ,\DSP_A_B_DATA.B2_DATA<12> ,\DSP_A_B_DATA.B2_DATA<11> ,\DSP_A_B_DATA.B2_DATA<10> ,\DSP_A_B_DATA.B2_DATA<9> ,\DSP_A_B_DATA.B2_DATA<8> ,\DSP_A_B_DATA.B2_DATA<7> ,\DSP_A_B_DATA.B2_DATA<6> ,\DSP_A_B_DATA.B2_DATA<5> ,\DSP_A_B_DATA.B2_DATA<4> ,\DSP_A_B_DATA.B2_DATA<3> ,\DSP_A_B_DATA.B2_DATA<2> ,\DSP_A_B_DATA.B2_DATA<1> ,\DSP_A_B_DATA.B2_DATA<0> }),
        .CEAD(CEAD),
        .CED(CED),
        .CEINMODE(CEINMODE),
        .CLK(CLK),
        .DIN({\D[26] ,\D[25] ,\D[24] ,\D[23] ,\D[22] ,\D[21] ,\D[20] ,\D[19] ,\D[18] ,\D[17] ,\D[16] ,\D[15] ,\D[14] ,\D[13] ,\D[12] ,\D[11] ,\D[10] ,\D[9] ,\D[8] ,\D[7] ,\D[6] ,\D[5] ,\D[4] ,\D[3] ,\D[2] ,\D[1] ,\D[0] }),
        .D_DATA({\DSP_PREADD_DATA.D_DATA<26> ,\DSP_PREADD_DATA.D_DATA<25> ,\DSP_PREADD_DATA.D_DATA<24> ,\DSP_PREADD_DATA.D_DATA<23> ,\DSP_PREADD_DATA.D_DATA<22> ,\DSP_PREADD_DATA.D_DATA<21> ,\DSP_PREADD_DATA.D_DATA<20> ,\DSP_PREADD_DATA.D_DATA<19> ,\DSP_PREADD_DATA.D_DATA<18> ,\DSP_PREADD_DATA.D_DATA<17> ,\DSP_PREADD_DATA.D_DATA<16> ,\DSP_PREADD_DATA.D_DATA<15> ,\DSP_PREADD_DATA.D_DATA<14> ,\DSP_PREADD_DATA.D_DATA<13> ,\DSP_PREADD_DATA.D_DATA<12> ,\DSP_PREADD_DATA.D_DATA<11> ,\DSP_PREADD_DATA.D_DATA<10> ,\DSP_PREADD_DATA.D_DATA<9> ,\DSP_PREADD_DATA.D_DATA<8> ,\DSP_PREADD_DATA.D_DATA<7> ,\DSP_PREADD_DATA.D_DATA<6> ,\DSP_PREADD_DATA.D_DATA<5> ,\DSP_PREADD_DATA.D_DATA<4> ,\DSP_PREADD_DATA.D_DATA<3> ,\DSP_PREADD_DATA.D_DATA<2> ,\DSP_PREADD_DATA.D_DATA<1> ,\DSP_PREADD_DATA.D_DATA<0> }),
        .INMODE({\INMODE[4] ,\INMODE[3] ,\INMODE[2] ,\INMODE[1] ,\INMODE[0] }),
        .INMODE_2(\DSP_PREADD_DATA.INMODE_2 ),
        .PREADD_AB({\DSP_PREADD_DATA.PREADD_AB<26> ,\DSP_PREADD_DATA.PREADD_AB<25> ,\DSP_PREADD_DATA.PREADD_AB<24> ,\DSP_PREADD_DATA.PREADD_AB<23> ,\DSP_PREADD_DATA.PREADD_AB<22> ,\DSP_PREADD_DATA.PREADD_AB<21> ,\DSP_PREADD_DATA.PREADD_AB<20> ,\DSP_PREADD_DATA.PREADD_AB<19> ,\DSP_PREADD_DATA.PREADD_AB<18> ,\DSP_PREADD_DATA.PREADD_AB<17> ,\DSP_PREADD_DATA.PREADD_AB<16> ,\DSP_PREADD_DATA.PREADD_AB<15> ,\DSP_PREADD_DATA.PREADD_AB<14> ,\DSP_PREADD_DATA.PREADD_AB<13> ,\DSP_PREADD_DATA.PREADD_AB<12> ,\DSP_PREADD_DATA.PREADD_AB<11> ,\DSP_PREADD_DATA.PREADD_AB<10> ,\DSP_PREADD_DATA.PREADD_AB<9> ,\DSP_PREADD_DATA.PREADD_AB<8> ,\DSP_PREADD_DATA.PREADD_AB<7> ,\DSP_PREADD_DATA.PREADD_AB<6> ,\DSP_PREADD_DATA.PREADD_AB<5> ,\DSP_PREADD_DATA.PREADD_AB<4> ,\DSP_PREADD_DATA.PREADD_AB<3> ,\DSP_PREADD_DATA.PREADD_AB<2> ,\DSP_PREADD_DATA.PREADD_AB<1> ,\DSP_PREADD_DATA.PREADD_AB<0> }),
        .RSTD(RSTD),
        .RSTINMODE(RSTINMODE));
  DSP_PREADD DSP_PREADD_INST
       (.AD({\DSP_PREADD.AD<26> ,\DSP_PREADD.AD<25> ,\DSP_PREADD.AD<24> ,\DSP_PREADD.AD<23> ,\DSP_PREADD.AD<22> ,\DSP_PREADD.AD<21> ,\DSP_PREADD.AD<20> ,\DSP_PREADD.AD<19> ,\DSP_PREADD.AD<18> ,\DSP_PREADD.AD<17> ,\DSP_PREADD.AD<16> ,\DSP_PREADD.AD<15> ,\DSP_PREADD.AD<14> ,\DSP_PREADD.AD<13> ,\DSP_PREADD.AD<12> ,\DSP_PREADD.AD<11> ,\DSP_PREADD.AD<10> ,\DSP_PREADD.AD<9> ,\DSP_PREADD.AD<8> ,\DSP_PREADD.AD<7> ,\DSP_PREADD.AD<6> ,\DSP_PREADD.AD<5> ,\DSP_PREADD.AD<4> ,\DSP_PREADD.AD<3> ,\DSP_PREADD.AD<2> ,\DSP_PREADD.AD<1> ,\DSP_PREADD.AD<0> }),
        .ADDSUB(\DSP_PREADD_DATA.ADDSUB ),
        .D_DATA({\DSP_PREADD_DATA.D_DATA<26> ,\DSP_PREADD_DATA.D_DATA<25> ,\DSP_PREADD_DATA.D_DATA<24> ,\DSP_PREADD_DATA.D_DATA<23> ,\DSP_PREADD_DATA.D_DATA<22> ,\DSP_PREADD_DATA.D_DATA<21> ,\DSP_PREADD_DATA.D_DATA<20> ,\DSP_PREADD_DATA.D_DATA<19> ,\DSP_PREADD_DATA.D_DATA<18> ,\DSP_PREADD_DATA.D_DATA<17> ,\DSP_PREADD_DATA.D_DATA<16> ,\DSP_PREADD_DATA.D_DATA<15> ,\DSP_PREADD_DATA.D_DATA<14> ,\DSP_PREADD_DATA.D_DATA<13> ,\DSP_PREADD_DATA.D_DATA<12> ,\DSP_PREADD_DATA.D_DATA<11> ,\DSP_PREADD_DATA.D_DATA<10> ,\DSP_PREADD_DATA.D_DATA<9> ,\DSP_PREADD_DATA.D_DATA<8> ,\DSP_PREADD_DATA.D_DATA<7> ,\DSP_PREADD_DATA.D_DATA<6> ,\DSP_PREADD_DATA.D_DATA<5> ,\DSP_PREADD_DATA.D_DATA<4> ,\DSP_PREADD_DATA.D_DATA<3> ,\DSP_PREADD_DATA.D_DATA<2> ,\DSP_PREADD_DATA.D_DATA<1> ,\DSP_PREADD_DATA.D_DATA<0> }),
        .INMODE2(\DSP_PREADD_DATA.INMODE_2 ),
        .PREADD_AB({\DSP_PREADD_DATA.PREADD_AB<26> ,\DSP_PREADD_DATA.PREADD_AB<25> ,\DSP_PREADD_DATA.PREADD_AB<24> ,\DSP_PREADD_DATA.PREADD_AB<23> ,\DSP_PREADD_DATA.PREADD_AB<22> ,\DSP_PREADD_DATA.PREADD_AB<21> ,\DSP_PREADD_DATA.PREADD_AB<20> ,\DSP_PREADD_DATA.PREADD_AB<19> ,\DSP_PREADD_DATA.PREADD_AB<18> ,\DSP_PREADD_DATA.PREADD_AB<17> ,\DSP_PREADD_DATA.PREADD_AB<16> ,\DSP_PREADD_DATA.PREADD_AB<15> ,\DSP_PREADD_DATA.PREADD_AB<14> ,\DSP_PREADD_DATA.PREADD_AB<13> ,\DSP_PREADD_DATA.PREADD_AB<12> ,\DSP_PREADD_DATA.PREADD_AB<11> ,\DSP_PREADD_DATA.PREADD_AB<10> ,\DSP_PREADD_DATA.PREADD_AB<9> ,\DSP_PREADD_DATA.PREADD_AB<8> ,\DSP_PREADD_DATA.PREADD_AB<7> ,\DSP_PREADD_DATA.PREADD_AB<6> ,\DSP_PREADD_DATA.PREADD_AB<5> ,\DSP_PREADD_DATA.PREADD_AB<4> ,\DSP_PREADD_DATA.PREADD_AB<3> ,\DSP_PREADD_DATA.PREADD_AB<2> ,\DSP_PREADD_DATA.PREADD_AB<1> ,\DSP_PREADD_DATA.PREADD_AB<0> }));
endmodule

module RAM32M16_UNIQ_BASE_
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32711
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32734
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32735
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32736
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32737
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32738
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM32M16_HD32739
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output [1:0]DOA;
  output [1:0]DOB;
  output [1:0]DOC;
  output [1:0]DOD;
  output [1:0]DOE;
  output [1:0]DOF;
  output [1:0]DOG;
  output [1:0]DOH;
  input [4:0]ADDRA;
  input [4:0]ADDRB;
  input [4:0]ADDRC;
  input [4:0]ADDRD;
  input [4:0]ADDRE;
  input [4:0]ADDRF;
  input [4:0]ADDRG;
  input [4:0]ADDRH;
  input [1:0]DIA;
  input [1:0]DIB;
  input [1:0]DIC;
  input [1:0]DID;
  input [1:0]DIE;
  input [1:0]DIF;
  input [1:0]DIG;
  input [1:0]DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire DIA0;
  wire DIA1;
  wire DIB0;
  wire DIB1;
  wire DIC0;
  wire DIC1;
  wire DID0;
  wire DID1;
  wire DIE0;
  wire DIE1;
  wire DIF0;
  wire DIF1;
  wire DIG0;
  wire DIG1;
  wire DIH0;
  wire DIH1;
  wire DOA0;
  wire DOA1;
  wire DOB0;
  wire DOB1;
  wire DOC0;
  wire DOC1;
  wire DOD0;
  wire DOD1;
  wire DOE0;
  wire DOE1;
  wire DOF0;
  wire DOF1;
  wire DOG0;
  wire DOG1;
  wire DOH0;
  wire DOH1;
  wire WCLK;
  wire WE;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign DIA0 = DIA[0];
  assign DIA1 = DIA[1];
  assign DIB0 = DIB[0];
  assign DIB1 = DIB[1];
  assign DIC0 = DIC[0];
  assign DIC1 = DIC[1];
  assign DID0 = DID[0];
  assign DID1 = DID[1];
  assign DIE0 = DIE[0];
  assign DIE1 = DIE[1];
  assign DIF0 = DIF[0];
  assign DIF1 = DIF[1];
  assign DIG0 = DIG[0];
  assign DIG1 = DIG[1];
  assign DIH0 = DIH[0];
  assign DIH1 = DIH[1];
  assign DOA[1] = DOA1;
  assign DOA[0] = DOA0;
  assign DOB[1] = DOB1;
  assign DOB[0] = DOB0;
  assign DOC[1] = DOC1;
  assign DOC[0] = DOC0;
  assign DOD[1] = DOD1;
  assign DOD[0] = DOD0;
  assign DOE[1] = DOE1;
  assign DOE[0] = DOE0;
  assign DOF[1] = DOF1;
  assign DOF[0] = DOF0;
  assign DOG[1] = DOG1;
  assign DOG[0] = DOG0;
  assign DOH[1] = DOH1;
  assign DOH[0] = DOH0;
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA0),
        .O(DOA0),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMA_D1
       (.CLK(WCLK),
        .I(DIA1),
        .O(DOA1),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB0),
        .O(DOB0),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMB_D1
       (.CLK(WCLK),
        .I(DIB1),
        .O(DOB1),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC0),
        .O(DOC0),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMC_D1
       (.CLK(WCLK),
        .I(DIC1),
        .O(DOC1),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD
       (.CLK(WCLK),
        .I(DID0),
        .O(DOD0),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMD_D1
       (.CLK(WCLK),
        .I(DID1),
        .O(DOD1),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME
       (.CLK(WCLK),
        .I(DIE0),
        .O(DOE0),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAME_D1
       (.CLK(WCLK),
        .I(DIE1),
        .O(DOE1),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF0),
        .O(DOF0),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMF_D1
       (.CLK(WCLK),
        .I(DIF1),
        .O(DOF1),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG0),
        .O(DOG0),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMD32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMG_D1
       (.CLK(WCLK),
        .I(DIG1),
        .O(DOG1),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH0),
        .O(DOH0),
        .WE(WE));
  RAMS32 #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    RAMH_D1
       (.ADR0(ADDRH0),
        .ADR1(ADDRH1),
        .ADR2(ADDRH2),
        .ADR3(ADDRH3),
        .ADR4(ADDRH4),
        .CLK(WCLK),
        .I(DIH1),
        .O(DOH1),
        .WE(WE));
endmodule

module RAM64M8_UNIQ_BASE_
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32712
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32714
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32715
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32716
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32717
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32718
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32719
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32720
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32721
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32723
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32724
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32725
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32726
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32727
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32728
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32729
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32730
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32731
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD32733
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64X1D_UNIQ_BASE_
   (DPO,
    SPO,
    A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    D,
    DPRA0,
    DPRA1,
    DPRA2,
    DPRA3,
    DPRA4,
    DPRA5,
    WCLK,
    WE);
  output DPO;
  output SPO;
  input A0;
  input A1;
  input A2;
  input A3;
  input A4;
  input A5;
  input D;
  input DPRA0;
  input DPRA1;
  input DPRA2;
  input DPRA3;
  input DPRA4;
  input DPRA5;
  input WCLK;
  input WE;

  wire A0;
  wire A1;
  wire A2;
  wire A3;
  wire A4;
  wire A5;
  wire D;
  wire DPO;
  wire DPRA0;
  wire DPRA1;
  wire DPRA2;
  wire DPRA3;
  wire DPRA4;
  wire DPRA5;
  wire SPO;
  wire WCLK;
  wire WE;
  wire NLW_DP_WADR6_UNCONNECTED;
  wire NLW_DP_WADR7_UNCONNECTED;
  wire NLW_SP_WADR6_UNCONNECTED;
  wire NLW_SP_WADR7_UNCONNECTED;

  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    DP
       (.CLK(WCLK),
        .I(D),
        .O(DPO),
        .RADR0(DPRA0),
        .RADR1(DPRA1),
        .RADR2(DPRA2),
        .RADR3(DPRA3),
        .RADR4(DPRA4),
        .RADR5(DPRA5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_DP_WADR6_UNCONNECTED),
        .WADR7(NLW_DP_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    SP
       (.CLK(WCLK),
        .I(D),
        .O(SPO),
        .RADR0(A0),
        .RADR1(A1),
        .RADR2(A2),
        .RADR3(A3),
        .RADR4(A4),
        .RADR5(A5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_SP_WADR6_UNCONNECTED),
        .WADR7(NLW_SP_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64X1D_HD32713
   (DPO,
    SPO,
    A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    D,
    DPRA0,
    DPRA1,
    DPRA2,
    DPRA3,
    DPRA4,
    DPRA5,
    WCLK,
    WE);
  output DPO;
  output SPO;
  input A0;
  input A1;
  input A2;
  input A3;
  input A4;
  input A5;
  input D;
  input DPRA0;
  input DPRA1;
  input DPRA2;
  input DPRA3;
  input DPRA4;
  input DPRA5;
  input WCLK;
  input WE;

  wire A0;
  wire A1;
  wire A2;
  wire A3;
  wire A4;
  wire A5;
  wire D;
  wire DPO;
  wire DPRA0;
  wire DPRA1;
  wire DPRA2;
  wire DPRA3;
  wire DPRA4;
  wire DPRA5;
  wire SPO;
  wire WCLK;
  wire WE;
  wire NLW_DP_WADR6_UNCONNECTED;
  wire NLW_DP_WADR7_UNCONNECTED;
  wire NLW_SP_WADR6_UNCONNECTED;
  wire NLW_SP_WADR7_UNCONNECTED;

  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    DP
       (.CLK(WCLK),
        .I(D),
        .O(DPO),
        .RADR0(DPRA0),
        .RADR1(DPRA1),
        .RADR2(DPRA2),
        .RADR3(DPRA3),
        .RADR4(DPRA4),
        .RADR5(DPRA5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_DP_WADR6_UNCONNECTED),
        .WADR7(NLW_DP_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    SP
       (.CLK(WCLK),
        .I(D),
        .O(SPO),
        .RADR0(A0),
        .RADR1(A1),
        .RADR2(A2),
        .RADR3(A3),
        .RADR4(A4),
        .RADR5(A5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_SP_WADR6_UNCONNECTED),
        .WADR7(NLW_SP_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64X1D_HD32722
   (DPO,
    SPO,
    A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    D,
    DPRA0,
    DPRA1,
    DPRA2,
    DPRA3,
    DPRA4,
    DPRA5,
    WCLK,
    WE);
  output DPO;
  output SPO;
  input A0;
  input A1;
  input A2;
  input A3;
  input A4;
  input A5;
  input D;
  input DPRA0;
  input DPRA1;
  input DPRA2;
  input DPRA3;
  input DPRA4;
  input DPRA5;
  input WCLK;
  input WE;

  wire A0;
  wire A1;
  wire A2;
  wire A3;
  wire A4;
  wire A5;
  wire D;
  wire DPO;
  wire DPRA0;
  wire DPRA1;
  wire DPRA2;
  wire DPRA3;
  wire DPRA4;
  wire DPRA5;
  wire SPO;
  wire WCLK;
  wire WE;
  wire NLW_DP_WADR6_UNCONNECTED;
  wire NLW_DP_WADR7_UNCONNECTED;
  wire NLW_SP_WADR6_UNCONNECTED;
  wire NLW_SP_WADR7_UNCONNECTED;

  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    DP
       (.CLK(WCLK),
        .I(D),
        .O(DPO),
        .RADR0(DPRA0),
        .RADR1(DPRA1),
        .RADR2(DPRA2),
        .RADR3(DPRA3),
        .RADR4(DPRA4),
        .RADR5(DPRA5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_DP_WADR6_UNCONNECTED),
        .WADR7(NLW_DP_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    SP
       (.CLK(WCLK),
        .I(D),
        .O(SPO),
        .RADR0(A0),
        .RADR1(A1),
        .RADR2(A2),
        .RADR3(A3),
        .RADR4(A4),
        .RADR5(A5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_SP_WADR6_UNCONNECTED),
        .WADR7(NLW_SP_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64X1D_HD32732
   (DPO,
    SPO,
    A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    D,
    DPRA0,
    DPRA1,
    DPRA2,
    DPRA3,
    DPRA4,
    DPRA5,
    WCLK,
    WE);
  output DPO;
  output SPO;
  input A0;
  input A1;
  input A2;
  input A3;
  input A4;
  input A5;
  input D;
  input DPRA0;
  input DPRA1;
  input DPRA2;
  input DPRA3;
  input DPRA4;
  input DPRA5;
  input WCLK;
  input WE;

  wire A0;
  wire A1;
  wire A2;
  wire A3;
  wire A4;
  wire A5;
  wire D;
  wire DPO;
  wire DPRA0;
  wire DPRA1;
  wire DPRA2;
  wire DPRA3;
  wire DPRA4;
  wire DPRA5;
  wire SPO;
  wire WCLK;
  wire WE;
  wire NLW_DP_WADR6_UNCONNECTED;
  wire NLW_DP_WADR7_UNCONNECTED;
  wire NLW_SP_WADR6_UNCONNECTED;
  wire NLW_SP_WADR7_UNCONNECTED;

  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    DP
       (.CLK(WCLK),
        .I(D),
        .O(DPO),
        .RADR0(DPRA0),
        .RADR1(DPRA1),
        .RADR2(DPRA2),
        .RADR3(DPRA3),
        .RADR4(DPRA4),
        .RADR5(DPRA5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_DP_WADR6_UNCONNECTED),
        .WADR7(NLW_DP_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    SP
       (.CLK(WCLK),
        .I(D),
        .O(SPO),
        .RADR0(A0),
        .RADR1(A1),
        .RADR2(A2),
        .RADR3(A3),
        .RADR4(A4),
        .RADR5(A5),
        .WADR0(A0),
        .WADR1(A1),
        .WADR2(A2),
        .WADR3(A3),
        .WADR4(A4),
        .WADR5(A5),
        .WADR6(NLW_SP_WADR6_UNCONNECTED),
        .WADR7(NLW_SP_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

(* dont_touch = "true" *) 
(* NotValidForBitStream *)
module switch_elements
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  (* DONT_TOUCH *) wire [15:0]DI;
  wire \DI_reg[15]_i_1_n_2 ;
  wire \DI_reg[15]_i_1_n_3 ;
  wire \DI_reg[15]_i_1_n_4 ;
  wire \DI_reg[15]_i_1_n_5 ;
  wire \DI_reg[15]_i_1_n_6 ;
  wire \DI_reg[15]_i_1_n_7 ;
  wire \DI_reg[8]_i_1_n_0 ;
  wire \DI_reg[8]_i_1_n_1 ;
  wire \DI_reg[8]_i_1_n_2 ;
  wire \DI_reg[8]_i_1_n_3 ;
  wire \DI_reg[8]_i_1_n_4 ;
  wire \DI_reg[8]_i_1_n_5 ;
  wire \DI_reg[8]_i_1_n_6 ;
  wire \DI_reg[8]_i_1_n_7 ;
  (* DONT_TOUCH *) wire [15:0]DO;
  (* DONT_TOUCH *) wire EF;
  (* DONT_TOUCH *) wire [15:0]FC_TRANS_PAUSEDATA;
  wire \FC_TRANS_PAUSEDATA[0]_i_1_n_0 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_10 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_11 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_12 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_13 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_14 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_15 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_2 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_3 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_4 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_5 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_6 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_7 ;
  wire \FC_TRANS_PAUSEDATA_reg[15]_i_1_n_9 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_0 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_1 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_10 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_11 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_12 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_13 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_14 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_15 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_2 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_3 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_4 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_5 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_6 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_7 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_8 ;
  wire \FC_TRANS_PAUSEDATA_reg[8]_i_1_n_9 ;
  (* DONT_TOUCH *) wire FC_TRANS_PAUSEVAL;
  (* DONT_TOUCH *) wire [15:0]FC_TX_PAUSEDATA;
  wire \FC_TX_PAUSEDATA[0]_i_1_n_0 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_10 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_11 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_12 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_13 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_14 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_15 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_2 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_3 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_4 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_5 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_6 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_7 ;
  wire \FC_TX_PAUSEDATA_reg[15]_i_1_n_9 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_0 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_1 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_10 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_11 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_12 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_13 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_14 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_15 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_2 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_3 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_4 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_5 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_6 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_7 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_8 ;
  wire \FC_TX_PAUSEDATA_reg[8]_i_1_n_9 ;
  (* DONT_TOUCH *) wire FC_TX_PAUSEVALID;
  (* DONT_TOUCH *) wire [11:0]FREQ;
  (* DONT_TOUCH *) wire LOCALLINKFAULT;
  (* DONT_TOUCH *) wire RXTXLINKFAULT;
  (* DONT_TOUCH *) wire [7:0]TXC;
  (* DONT_TOUCH *) wire [63:0]TXD;
  (* DONT_TOUCH *) wire TX_ACK;
  (* DONT_TOUCH *) wire TX_CFG_REG_VALID;
  (* DONT_TOUCH *) wire [31:0]TX_CFG_REG_VALUE;
  (* DONT_TOUCH *) wire [63:0]TX_DATA;
  wire \TX_DATA[0]_i_1_n_0 ;
  (* DONT_TOUCH *) wire [7:0]TX_DATA_VALID;
  wire \TX_DATA_VALID[0]_i_1_n_0 ;
  wire \TX_DATA_VALID[1]_i_1_n_0 ;
  wire \TX_DATA_VALID[2]_i_1_n_0 ;
  wire \TX_DATA_VALID[3]_i_1_n_0 ;
  wire \TX_DATA_VALID[4]_i_1_n_0 ;
  wire \TX_DATA_VALID[5]_i_1_n_0 ;
  wire \TX_DATA_VALID[6]_i_1_n_0 ;
  wire \TX_DATA_VALID[7]_i_1_n_0 ;
  wire \TX_DATA_VALID[7]_i_2_n_0 ;
  wire \TX_DATA_reg[16]_i_1_n_0 ;
  wire \TX_DATA_reg[16]_i_1_n_1 ;
  wire \TX_DATA_reg[16]_i_1_n_10 ;
  wire \TX_DATA_reg[16]_i_1_n_11 ;
  wire \TX_DATA_reg[16]_i_1_n_12 ;
  wire \TX_DATA_reg[16]_i_1_n_13 ;
  wire \TX_DATA_reg[16]_i_1_n_14 ;
  wire \TX_DATA_reg[16]_i_1_n_15 ;
  wire \TX_DATA_reg[16]_i_1_n_2 ;
  wire \TX_DATA_reg[16]_i_1_n_3 ;
  wire \TX_DATA_reg[16]_i_1_n_4 ;
  wire \TX_DATA_reg[16]_i_1_n_5 ;
  wire \TX_DATA_reg[16]_i_1_n_6 ;
  wire \TX_DATA_reg[16]_i_1_n_7 ;
  wire \TX_DATA_reg[16]_i_1_n_8 ;
  wire \TX_DATA_reg[16]_i_1_n_9 ;
  wire \TX_DATA_reg[24]_i_1_n_0 ;
  wire \TX_DATA_reg[24]_i_1_n_1 ;
  wire \TX_DATA_reg[24]_i_1_n_10 ;
  wire \TX_DATA_reg[24]_i_1_n_11 ;
  wire \TX_DATA_reg[24]_i_1_n_12 ;
  wire \TX_DATA_reg[24]_i_1_n_13 ;
  wire \TX_DATA_reg[24]_i_1_n_14 ;
  wire \TX_DATA_reg[24]_i_1_n_15 ;
  wire \TX_DATA_reg[24]_i_1_n_2 ;
  wire \TX_DATA_reg[24]_i_1_n_3 ;
  wire \TX_DATA_reg[24]_i_1_n_4 ;
  wire \TX_DATA_reg[24]_i_1_n_5 ;
  wire \TX_DATA_reg[24]_i_1_n_6 ;
  wire \TX_DATA_reg[24]_i_1_n_7 ;
  wire \TX_DATA_reg[24]_i_1_n_8 ;
  wire \TX_DATA_reg[24]_i_1_n_9 ;
  wire \TX_DATA_reg[32]_i_1_n_0 ;
  wire \TX_DATA_reg[32]_i_1_n_1 ;
  wire \TX_DATA_reg[32]_i_1_n_10 ;
  wire \TX_DATA_reg[32]_i_1_n_11 ;
  wire \TX_DATA_reg[32]_i_1_n_12 ;
  wire \TX_DATA_reg[32]_i_1_n_13 ;
  wire \TX_DATA_reg[32]_i_1_n_14 ;
  wire \TX_DATA_reg[32]_i_1_n_15 ;
  wire \TX_DATA_reg[32]_i_1_n_2 ;
  wire \TX_DATA_reg[32]_i_1_n_3 ;
  wire \TX_DATA_reg[32]_i_1_n_4 ;
  wire \TX_DATA_reg[32]_i_1_n_5 ;
  wire \TX_DATA_reg[32]_i_1_n_6 ;
  wire \TX_DATA_reg[32]_i_1_n_7 ;
  wire \TX_DATA_reg[32]_i_1_n_8 ;
  wire \TX_DATA_reg[32]_i_1_n_9 ;
  wire \TX_DATA_reg[40]_i_1_n_0 ;
  wire \TX_DATA_reg[40]_i_1_n_1 ;
  wire \TX_DATA_reg[40]_i_1_n_10 ;
  wire \TX_DATA_reg[40]_i_1_n_11 ;
  wire \TX_DATA_reg[40]_i_1_n_12 ;
  wire \TX_DATA_reg[40]_i_1_n_13 ;
  wire \TX_DATA_reg[40]_i_1_n_14 ;
  wire \TX_DATA_reg[40]_i_1_n_15 ;
  wire \TX_DATA_reg[40]_i_1_n_2 ;
  wire \TX_DATA_reg[40]_i_1_n_3 ;
  wire \TX_DATA_reg[40]_i_1_n_4 ;
  wire \TX_DATA_reg[40]_i_1_n_5 ;
  wire \TX_DATA_reg[40]_i_1_n_6 ;
  wire \TX_DATA_reg[40]_i_1_n_7 ;
  wire \TX_DATA_reg[40]_i_1_n_8 ;
  wire \TX_DATA_reg[40]_i_1_n_9 ;
  wire \TX_DATA_reg[48]_i_1_n_0 ;
  wire \TX_DATA_reg[48]_i_1_n_1 ;
  wire \TX_DATA_reg[48]_i_1_n_10 ;
  wire \TX_DATA_reg[48]_i_1_n_11 ;
  wire \TX_DATA_reg[48]_i_1_n_12 ;
  wire \TX_DATA_reg[48]_i_1_n_13 ;
  wire \TX_DATA_reg[48]_i_1_n_14 ;
  wire \TX_DATA_reg[48]_i_1_n_15 ;
  wire \TX_DATA_reg[48]_i_1_n_2 ;
  wire \TX_DATA_reg[48]_i_1_n_3 ;
  wire \TX_DATA_reg[48]_i_1_n_4 ;
  wire \TX_DATA_reg[48]_i_1_n_5 ;
  wire \TX_DATA_reg[48]_i_1_n_6 ;
  wire \TX_DATA_reg[48]_i_1_n_7 ;
  wire \TX_DATA_reg[48]_i_1_n_8 ;
  wire \TX_DATA_reg[48]_i_1_n_9 ;
  wire \TX_DATA_reg[56]_i_1_n_0 ;
  wire \TX_DATA_reg[56]_i_1_n_1 ;
  wire \TX_DATA_reg[56]_i_1_n_10 ;
  wire \TX_DATA_reg[56]_i_1_n_11 ;
  wire \TX_DATA_reg[56]_i_1_n_12 ;
  wire \TX_DATA_reg[56]_i_1_n_13 ;
  wire \TX_DATA_reg[56]_i_1_n_14 ;
  wire \TX_DATA_reg[56]_i_1_n_15 ;
  wire \TX_DATA_reg[56]_i_1_n_2 ;
  wire \TX_DATA_reg[56]_i_1_n_3 ;
  wire \TX_DATA_reg[56]_i_1_n_4 ;
  wire \TX_DATA_reg[56]_i_1_n_5 ;
  wire \TX_DATA_reg[56]_i_1_n_6 ;
  wire \TX_DATA_reg[56]_i_1_n_7 ;
  wire \TX_DATA_reg[56]_i_1_n_8 ;
  wire \TX_DATA_reg[56]_i_1_n_9 ;
  wire \TX_DATA_reg[63]_i_1_n_10 ;
  wire \TX_DATA_reg[63]_i_1_n_11 ;
  wire \TX_DATA_reg[63]_i_1_n_12 ;
  wire \TX_DATA_reg[63]_i_1_n_13 ;
  wire \TX_DATA_reg[63]_i_1_n_14 ;
  wire \TX_DATA_reg[63]_i_1_n_15 ;
  wire \TX_DATA_reg[63]_i_1_n_2 ;
  wire \TX_DATA_reg[63]_i_1_n_3 ;
  wire \TX_DATA_reg[63]_i_1_n_4 ;
  wire \TX_DATA_reg[63]_i_1_n_5 ;
  wire \TX_DATA_reg[63]_i_1_n_6 ;
  wire \TX_DATA_reg[63]_i_1_n_7 ;
  wire \TX_DATA_reg[63]_i_1_n_9 ;
  wire \TX_DATA_reg[8]_i_1_n_0 ;
  wire \TX_DATA_reg[8]_i_1_n_1 ;
  wire \TX_DATA_reg[8]_i_1_n_10 ;
  wire \TX_DATA_reg[8]_i_1_n_11 ;
  wire \TX_DATA_reg[8]_i_1_n_12 ;
  wire \TX_DATA_reg[8]_i_1_n_13 ;
  wire \TX_DATA_reg[8]_i_1_n_14 ;
  wire \TX_DATA_reg[8]_i_1_n_15 ;
  wire \TX_DATA_reg[8]_i_1_n_2 ;
  wire \TX_DATA_reg[8]_i_1_n_3 ;
  wire \TX_DATA_reg[8]_i_1_n_4 ;
  wire \TX_DATA_reg[8]_i_1_n_5 ;
  wire \TX_DATA_reg[8]_i_1_n_6 ;
  wire \TX_DATA_reg[8]_i_1_n_7 ;
  wire \TX_DATA_reg[8]_i_1_n_8 ;
  wire \TX_DATA_reg[8]_i_1_n_9 ;
  (* DONT_TOUCH *) wire [7:0]TX_IFG_DELAY;
  wire \TX_IFG_DELAY[0]_i_1_n_0 ;
  wire \TX_IFG_DELAY[1]_i_1_n_0 ;
  wire \TX_IFG_DELAY[2]_i_1_n_0 ;
  wire \TX_IFG_DELAY[3]_i_1_n_0 ;
  wire \TX_IFG_DELAY[4]_i_1_n_0 ;
  wire \TX_IFG_DELAY[5]_i_1_n_0 ;
  wire \TX_IFG_DELAY[6]_i_1_n_0 ;
  wire \TX_IFG_DELAY[7]_i_1_n_0 ;
  wire \TX_IFG_DELAY[7]_i_2_n_0 ;
  (* DONT_TOUCH *) wire TX_START;
  (* DONT_TOUCH *) wire TX_STATS_VALID;
  (* DONT_TOUCH *) wire TX_UNDERRUN;
  (* DONT_TOUCH *) wire ack_o;
  wire \activity_blocks[0].dutH_n_0 ;
  wire activity_blocks_c_0_n_0;
  wire activity_blocks_c_10_n_0;
  wire activity_blocks_c_11_n_0;
  wire activity_blocks_c_1_n_0;
  wire activity_blocks_c_2_n_0;
  wire activity_blocks_c_3_n_0;
  wire activity_blocks_c_4_n_0;
  wire activity_blocks_c_5_n_0;
  wire activity_blocks_c_6_n_0;
  wire activity_blocks_c_7_n_0;
  wire activity_blocks_c_8_n_0;
  wire activity_blocks_c_9_n_0;
  wire activity_blocks_c_n_0;
  (* DONT_TOUCH *) wire [10:0]addr;
  wire \addr[0]_i_1_n_0 ;
  wire \addr[10]_i_1_n_0 ;
  wire \addr[10]_i_2_n_0 ;
  wire \addr[1]_i_1_n_0 ;
  wire \addr[2]_i_1_n_0 ;
  wire \addr[3]_i_1_n_0 ;
  wire \addr[4]_i_1_n_0 ;
  wire \addr[5]_i_1_n_0 ;
  wire \addr[6]_i_1_n_0 ;
  wire \addr[7]_i_1_n_0 ;
  wire \addr[8]_i_1_n_0 ;
  wire \addr[9]_i_1_n_0 ;
  (* DONT_TOUCH *) wire [1:0]adr_i;
  (* DONT_TOUCH *) wire [52:0]cfgRxRegData;
  (* DONT_TOUCH *) wire [64:0]cfgRxRegData_in;
  wire \cfgRxRegData_in[0]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[16]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[24]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[32]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[40]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[48]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[56]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[64]_i_1_n_9 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_0 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_1 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_10 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_11 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_12 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_13 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_14 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_15 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_2 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_3 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_4 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_5 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_6 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_7 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_8 ;
  wire \cfgRxRegData_in_reg[8]_i_1_n_9 ;
  (* DONT_TOUCH *) wire [9:0]cfgTxRegData;
  (* DONT_TOUCH *) wire crc_en;
  (* DONT_TOUCH *) wire cyc_i;
  wire d4_30;
  (* DONT_TOUCH *) wire dat_i;
  (* DONT_TOUCH *) wire [7:0]dat_i_vec;
  (* DONT_TOUCH *) wire [7:0]dat_o;
  (* DONT_TOUCH *) wire [4:0]dat_o_vec;
  (* DONT_TOUCH *) wire data_i;
  wire [31:0]info_o;
  wire \info_o[0]_INST_0_i_1_n_0 ;
  (* DONT_TOUCH *) wire [7:0]inputs;
  (* DONT_TOUCH *) wire inta_o;
  (* DONT_TOUCH *) wire m_en;
  (* DONT_TOUCH *) wire [1:0]m_we;
  (* DONT_TOUCH *) wire mdc;
  (* DONT_TOUCH *) wire mdio;
  (* DONT_TOUCH *) wire [9:0]mgmt_addr;
  (* DONT_TOUCH *) wire mgmt_miim_rdy;
  (* DONT_TOUCH *) wire mgmt_miim_sel;
  (* DONT_TOUCH *) wire [1:0]mgmt_opcode;
  (* DONT_TOUCH *) wire [31:0]mgmt_rd_data;
  (* DONT_TOUCH *) wire mgmt_req;
  (* DONT_TOUCH *) wire [31:0]mgmt_wr_data;
  (* DONT_TOUCH *) wire miso_i;
  (* DONT_TOUCH *) wire mosi_o;
  (* DONT_TOUCH *) wire [7:0]outputs;
  wire [15:0]plusOp;
  (* DONT_TOUCH *) wire [3:0]q_o;
  (* DONT_TOUCH *) wire [15:0]rdata;
  (* DONT_TOUCH *) wire ready_o;
  (* DONT_TOUCH *) wire [3:0]recieved_debug;
  wire rst_i;
  (* DONT_TOUCH *) wire rst_syn;
  (* DONT_TOUCH *) wire run_in;
  (* DONT_TOUCH *) wire run_out;
  (* DONT_TOUCH *) wire [2:0]rxCfgofRS;
  (* DONT_TOUCH *) wire [18:0]rxStatRegPlus;
  (* DONT_TOUCH *) wire [1:0]rxTxLinkFault_vec;
  (* DONT_TOUCH *) wire rx_bad_frame;
  (* DONT_TOUCH *) wire [63:0]rx_data;
  (* DONT_TOUCH *) wire [7:0]rx_data_valid;
  (* DONT_TOUCH *) wire rx_good_frame;
  wire rxclk_180;
  (* DONT_TOUCH *) wire rxclk_out;
  (* DONT_TOUCH *) wire sck_o;
  (* DONT_TOUCH *) wire stb_i;
  (* DONT_TOUCH *) wire [24:0]txStatRegPlus;
  (* DONT_TOUCH *) wire waitforstart_rdy;
  (* DONT_TOUCH *) wire [15:0]wdata;
  (* DONT_TOUCH *) wire we_i;
  (* DONT_TOUCH *) wire [3:0]xgmii_rxc;
  (* DONT_TOUCH *) wire [31:0]xgmii_rxd;
  wire \xgmii_rxd[0]_i_1_n_0 ;
  wire \xgmii_rxd_reg[16]_i_1_n_0 ;
  wire \xgmii_rxd_reg[16]_i_1_n_1 ;
  wire \xgmii_rxd_reg[16]_i_1_n_10 ;
  wire \xgmii_rxd_reg[16]_i_1_n_11 ;
  wire \xgmii_rxd_reg[16]_i_1_n_12 ;
  wire \xgmii_rxd_reg[16]_i_1_n_13 ;
  wire \xgmii_rxd_reg[16]_i_1_n_14 ;
  wire \xgmii_rxd_reg[16]_i_1_n_15 ;
  wire \xgmii_rxd_reg[16]_i_1_n_2 ;
  wire \xgmii_rxd_reg[16]_i_1_n_3 ;
  wire \xgmii_rxd_reg[16]_i_1_n_4 ;
  wire \xgmii_rxd_reg[16]_i_1_n_5 ;
  wire \xgmii_rxd_reg[16]_i_1_n_6 ;
  wire \xgmii_rxd_reg[16]_i_1_n_7 ;
  wire \xgmii_rxd_reg[16]_i_1_n_8 ;
  wire \xgmii_rxd_reg[16]_i_1_n_9 ;
  wire \xgmii_rxd_reg[24]_i_1_n_0 ;
  wire \xgmii_rxd_reg[24]_i_1_n_1 ;
  wire \xgmii_rxd_reg[24]_i_1_n_10 ;
  wire \xgmii_rxd_reg[24]_i_1_n_11 ;
  wire \xgmii_rxd_reg[24]_i_1_n_12 ;
  wire \xgmii_rxd_reg[24]_i_1_n_13 ;
  wire \xgmii_rxd_reg[24]_i_1_n_14 ;
  wire \xgmii_rxd_reg[24]_i_1_n_15 ;
  wire \xgmii_rxd_reg[24]_i_1_n_2 ;
  wire \xgmii_rxd_reg[24]_i_1_n_3 ;
  wire \xgmii_rxd_reg[24]_i_1_n_4 ;
  wire \xgmii_rxd_reg[24]_i_1_n_5 ;
  wire \xgmii_rxd_reg[24]_i_1_n_6 ;
  wire \xgmii_rxd_reg[24]_i_1_n_7 ;
  wire \xgmii_rxd_reg[24]_i_1_n_8 ;
  wire \xgmii_rxd_reg[24]_i_1_n_9 ;
  wire \xgmii_rxd_reg[31]_i_1_n_10 ;
  wire \xgmii_rxd_reg[31]_i_1_n_11 ;
  wire \xgmii_rxd_reg[31]_i_1_n_12 ;
  wire \xgmii_rxd_reg[31]_i_1_n_13 ;
  wire \xgmii_rxd_reg[31]_i_1_n_14 ;
  wire \xgmii_rxd_reg[31]_i_1_n_15 ;
  wire \xgmii_rxd_reg[31]_i_1_n_2 ;
  wire \xgmii_rxd_reg[31]_i_1_n_3 ;
  wire \xgmii_rxd_reg[31]_i_1_n_4 ;
  wire \xgmii_rxd_reg[31]_i_1_n_5 ;
  wire \xgmii_rxd_reg[31]_i_1_n_6 ;
  wire \xgmii_rxd_reg[31]_i_1_n_7 ;
  wire \xgmii_rxd_reg[31]_i_1_n_9 ;
  wire \xgmii_rxd_reg[8]_i_1_n_0 ;
  wire \xgmii_rxd_reg[8]_i_1_n_1 ;
  wire \xgmii_rxd_reg[8]_i_1_n_10 ;
  wire \xgmii_rxd_reg[8]_i_1_n_11 ;
  wire \xgmii_rxd_reg[8]_i_1_n_12 ;
  wire \xgmii_rxd_reg[8]_i_1_n_13 ;
  wire \xgmii_rxd_reg[8]_i_1_n_14 ;
  wire \xgmii_rxd_reg[8]_i_1_n_15 ;
  wire \xgmii_rxd_reg[8]_i_1_n_2 ;
  wire \xgmii_rxd_reg[8]_i_1_n_3 ;
  wire \xgmii_rxd_reg[8]_i_1_n_4 ;
  wire \xgmii_rxd_reg[8]_i_1_n_5 ;
  wire \xgmii_rxd_reg[8]_i_1_n_6 ;
  wire \xgmii_rxd_reg[8]_i_1_n_7 ;
  wire \xgmii_rxd_reg[8]_i_1_n_8 ;
  wire \xgmii_rxd_reg[8]_i_1_n_9 ;
  wire [7:6]\NLW_DI_reg[15]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_DI_reg[15]_i_1_O_UNCONNECTED ;
  wire [7:6]\NLW_FC_TRANS_PAUSEDATA_reg[15]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_FC_TRANS_PAUSEDATA_reg[15]_i_1_O_UNCONNECTED ;
  wire [7:6]\NLW_FC_TX_PAUSEDATA_reg[15]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_FC_TX_PAUSEDATA_reg[15]_i_1_O_UNCONNECTED ;
  wire [7:6]\NLW_TX_DATA_reg[63]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_TX_DATA_reg[63]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_cfgRxRegData_in_reg[64]_i_1_CO_UNCONNECTED ;
  wire [7:6]\NLW_xgmii_rxd_reg[31]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_xgmii_rxd_reg[31]_i_1_O_UNCONNECTED ;

  assign crc_en = enable_i[0];
  assign dat_i = enable_i[7];
  assign inputs = enable_i[31:24];
  assign mgmt_wr_data[23:16] = enable_i[23:16];
  assign rxclk_out = clk_i;
  assign wdata[15:8] = enable_i[15:8];
  assign wdata[6:1] = enable_i[6:1];
  LUT1 #(
    .INIT(2'h1)) 
    \DI[0]_i_1 
       (.I0(DI[0]),
        .O(plusOp[0]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[0]),
        .Q(DI[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[10]),
        .Q(DI[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[11] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[11]),
        .Q(DI[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[12] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[12]),
        .Q(DI[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[13] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[13]),
        .Q(DI[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[14] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[14]),
        .Q(DI[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[15] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[15]),
        .Q(DI[15]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \DI_reg[15]_i_1 
       (.CI(\DI_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_DI_reg[15]_i_1_CO_UNCONNECTED [7:6],\DI_reg[15]_i_1_n_2 ,\DI_reg[15]_i_1_n_3 ,\DI_reg[15]_i_1_n_4 ,\DI_reg[15]_i_1_n_5 ,\DI_reg[15]_i_1_n_6 ,\DI_reg[15]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_DI_reg[15]_i_1_O_UNCONNECTED [7],plusOp[15:9]}),
        .S({1'b0,DI[15:9]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[1]),
        .Q(DI[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[2]),
        .Q(DI[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[3]),
        .Q(DI[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[4]),
        .Q(DI[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[5]),
        .Q(DI[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[6]),
        .Q(DI[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[7]),
        .Q(DI[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[8]),
        .Q(DI[8]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \DI_reg[8]_i_1 
       (.CI(DI[0]),
        .CI_TOP(1'b0),
        .CO({\DI_reg[8]_i_1_n_0 ,\DI_reg[8]_i_1_n_1 ,\DI_reg[8]_i_1_n_2 ,\DI_reg[8]_i_1_n_3 ,\DI_reg[8]_i_1_n_4 ,\DI_reg[8]_i_1_n_5 ,\DI_reg[8]_i_1_n_6 ,\DI_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(plusOp[8:1]),
        .S(DI[8:1]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DI_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(plusOp[9]),
        .Q(DI[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h2)) 
    EF_inst
       (.I0(wdata[3]),
        .O(EF));
  LUT1 #(
    .INIT(2'h1)) 
    \FC_TRANS_PAUSEDATA[0]_i_1 
       (.I0(FC_TRANS_PAUSEDATA[0]),
        .O(\FC_TRANS_PAUSEDATA[0]_i_1_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA[0]_i_1_n_0 ),
        .Q(FC_TRANS_PAUSEDATA[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_14 ),
        .Q(FC_TRANS_PAUSEDATA[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[11] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_13 ),
        .Q(FC_TRANS_PAUSEDATA[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[12] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_12 ),
        .Q(FC_TRANS_PAUSEDATA[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[13] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_11 ),
        .Q(FC_TRANS_PAUSEDATA[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[14] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_10 ),
        .Q(FC_TRANS_PAUSEDATA[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[15] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_9 ),
        .Q(FC_TRANS_PAUSEDATA[15]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \FC_TRANS_PAUSEDATA_reg[15]_i_1 
       (.CI(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_FC_TRANS_PAUSEDATA_reg[15]_i_1_CO_UNCONNECTED [7:6],\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_2 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_3 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_4 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_5 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_6 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_FC_TRANS_PAUSEDATA_reg[15]_i_1_O_UNCONNECTED [7],\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_9 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_10 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_11 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_12 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_13 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_14 ,\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_15 }),
        .S({1'b0,FC_TRANS_PAUSEDATA[15:9]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_15 ),
        .Q(FC_TRANS_PAUSEDATA[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_14 ),
        .Q(FC_TRANS_PAUSEDATA[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_13 ),
        .Q(FC_TRANS_PAUSEDATA[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_12 ),
        .Q(FC_TRANS_PAUSEDATA[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_11 ),
        .Q(FC_TRANS_PAUSEDATA[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_10 ),
        .Q(FC_TRANS_PAUSEDATA[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_9 ),
        .Q(FC_TRANS_PAUSEDATA[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_8 ),
        .Q(FC_TRANS_PAUSEDATA[8]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \FC_TRANS_PAUSEDATA_reg[8]_i_1 
       (.CI(FC_TRANS_PAUSEDATA[0]),
        .CI_TOP(1'b0),
        .CO({\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_0 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_1 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_2 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_3 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_4 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_5 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_6 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_8 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_9 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_10 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_11 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_12 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_13 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_14 ,\FC_TRANS_PAUSEDATA_reg[8]_i_1_n_15 }),
        .S(FC_TRANS_PAUSEDATA[8:1]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TRANS_PAUSEDATA_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TRANS_PAUSEDATA_reg[15]_i_1_n_15 ),
        .Q(FC_TRANS_PAUSEDATA[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h2)) 
    FC_TRANS_PAUSEVAL_inst
       (.I0(wdata[1]),
        .O(FC_TRANS_PAUSEVAL));
  LUT1 #(
    .INIT(2'h1)) 
    \FC_TX_PAUSEDATA[0]_i_1 
       (.I0(FC_TX_PAUSEDATA[0]),
        .O(\FC_TX_PAUSEDATA[0]_i_1_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA[0]_i_1_n_0 ),
        .Q(FC_TX_PAUSEDATA[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_14 ),
        .Q(FC_TX_PAUSEDATA[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[11] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_13 ),
        .Q(FC_TX_PAUSEDATA[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[12] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_12 ),
        .Q(FC_TX_PAUSEDATA[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[13] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_11 ),
        .Q(FC_TX_PAUSEDATA[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[14] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_10 ),
        .Q(FC_TX_PAUSEDATA[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[15] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_9 ),
        .Q(FC_TX_PAUSEDATA[15]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \FC_TX_PAUSEDATA_reg[15]_i_1 
       (.CI(\FC_TX_PAUSEDATA_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_FC_TX_PAUSEDATA_reg[15]_i_1_CO_UNCONNECTED [7:6],\FC_TX_PAUSEDATA_reg[15]_i_1_n_2 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_3 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_4 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_5 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_6 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_FC_TX_PAUSEDATA_reg[15]_i_1_O_UNCONNECTED [7],\FC_TX_PAUSEDATA_reg[15]_i_1_n_9 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_10 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_11 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_12 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_13 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_14 ,\FC_TX_PAUSEDATA_reg[15]_i_1_n_15 }),
        .S({1'b0,FC_TX_PAUSEDATA[15:9]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_15 ),
        .Q(FC_TX_PAUSEDATA[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_14 ),
        .Q(FC_TX_PAUSEDATA[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_13 ),
        .Q(FC_TX_PAUSEDATA[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_12 ),
        .Q(FC_TX_PAUSEDATA[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_11 ),
        .Q(FC_TX_PAUSEDATA[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_10 ),
        .Q(FC_TX_PAUSEDATA[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_9 ),
        .Q(FC_TX_PAUSEDATA[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[8]_i_1_n_8 ),
        .Q(FC_TX_PAUSEDATA[8]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \FC_TX_PAUSEDATA_reg[8]_i_1 
       (.CI(FC_TX_PAUSEDATA[0]),
        .CI_TOP(1'b0),
        .CO({\FC_TX_PAUSEDATA_reg[8]_i_1_n_0 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_1 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_2 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_3 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_4 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_5 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_6 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\FC_TX_PAUSEDATA_reg[8]_i_1_n_8 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_9 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_10 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_11 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_12 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_13 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_14 ,\FC_TX_PAUSEDATA_reg[8]_i_1_n_15 }),
        .S(FC_TX_PAUSEDATA[8:1]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FC_TX_PAUSEDATA_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\FC_TX_PAUSEDATA_reg[15]_i_1_n_15 ),
        .Q(FC_TX_PAUSEDATA[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h2)) 
    FC_TX_PAUSEVALID_inst
       (.I0(wdata[2]),
        .O(FC_TX_PAUSEVALID));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst
       (.I0(inputs[3]),
        .O(FREQ[11]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__0
       (.I0(inputs[2]),
        .O(FREQ[10]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__1
       (.I0(inputs[1]),
        .O(FREQ[9]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__10
       (.I0(mgmt_wr_data[16]),
        .O(FREQ[0]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__2
       (.I0(inputs[0]),
        .O(FREQ[8]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__3
       (.I0(mgmt_wr_data[23]),
        .O(FREQ[7]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__4
       (.I0(mgmt_wr_data[22]),
        .O(FREQ[6]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__5
       (.I0(mgmt_wr_data[21]),
        .O(FREQ[5]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__6
       (.I0(mgmt_wr_data[20]),
        .O(FREQ[4]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__7
       (.I0(mgmt_wr_data[19]),
        .O(FREQ[3]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__8
       (.I0(mgmt_wr_data[18]),
        .O(FREQ[2]));
  LUT1 #(
    .INIT(2'h2)) 
    FREQ_inst__9
       (.I0(mgmt_wr_data[17]),
        .O(FREQ[1]));
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_linkstate_reg[1]_i_3 
       (.I0(rxclk_out),
        .O(rxclk_180));
  LUT1 #(
    .INIT(2'h2)) 
    LOCALLINKFAULT_inst
       (.I0(inputs[7]),
        .O(LOCALLINKFAULT));
  LUT1 #(
    .INIT(2'h2)) 
    RXTXLINKFAULT_inst
       (.I0(wdata[2]),
        .O(RXTXLINKFAULT));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALID_inst
       (.I0(crc_en),
        .O(TX_CFG_REG_VALID));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst
       (.I0(inputs[7]),
        .O(TX_CFG_REG_VALUE[31]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__0
       (.I0(inputs[6]),
        .O(TX_CFG_REG_VALUE[30]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__1
       (.I0(inputs[5]),
        .O(TX_CFG_REG_VALUE[29]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__10
       (.I0(mgmt_wr_data[20]),
        .O(TX_CFG_REG_VALUE[20]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__11
       (.I0(mgmt_wr_data[19]),
        .O(TX_CFG_REG_VALUE[19]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__12
       (.I0(mgmt_wr_data[18]),
        .O(TX_CFG_REG_VALUE[18]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__13
       (.I0(mgmt_wr_data[17]),
        .O(TX_CFG_REG_VALUE[17]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__14
       (.I0(mgmt_wr_data[16]),
        .O(TX_CFG_REG_VALUE[16]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__15
       (.I0(wdata[15]),
        .O(TX_CFG_REG_VALUE[15]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__16
       (.I0(wdata[14]),
        .O(TX_CFG_REG_VALUE[14]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__17
       (.I0(wdata[13]),
        .O(TX_CFG_REG_VALUE[13]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__18
       (.I0(wdata[12]),
        .O(TX_CFG_REG_VALUE[12]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__19
       (.I0(wdata[11]),
        .O(TX_CFG_REG_VALUE[11]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__2
       (.I0(inputs[4]),
        .O(TX_CFG_REG_VALUE[28]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__20
       (.I0(wdata[10]),
        .O(TX_CFG_REG_VALUE[10]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__21
       (.I0(wdata[9]),
        .O(TX_CFG_REG_VALUE[9]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__22
       (.I0(wdata[8]),
        .O(TX_CFG_REG_VALUE[8]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__23
       (.I0(dat_i),
        .O(TX_CFG_REG_VALUE[7]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__24
       (.I0(wdata[6]),
        .O(TX_CFG_REG_VALUE[6]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__25
       (.I0(wdata[5]),
        .O(TX_CFG_REG_VALUE[5]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__26
       (.I0(wdata[4]),
        .O(TX_CFG_REG_VALUE[4]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__27
       (.I0(wdata[3]),
        .O(TX_CFG_REG_VALUE[3]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__28
       (.I0(wdata[2]),
        .O(TX_CFG_REG_VALUE[2]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__29
       (.I0(wdata[1]),
        .O(TX_CFG_REG_VALUE[1]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__3
       (.I0(inputs[3]),
        .O(TX_CFG_REG_VALUE[27]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__30
       (.I0(crc_en),
        .O(TX_CFG_REG_VALUE[0]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__4
       (.I0(inputs[2]),
        .O(TX_CFG_REG_VALUE[26]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__5
       (.I0(inputs[1]),
        .O(TX_CFG_REG_VALUE[25]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__6
       (.I0(inputs[0]),
        .O(TX_CFG_REG_VALUE[24]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__7
       (.I0(mgmt_wr_data[23]),
        .O(TX_CFG_REG_VALUE[23]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__8
       (.I0(mgmt_wr_data[22]),
        .O(TX_CFG_REG_VALUE[22]));
  LUT1 #(
    .INIT(2'h2)) 
    TX_CFG_REG_VALUE_inst__9
       (.I0(mgmt_wr_data[21]),
        .O(TX_CFG_REG_VALUE[21]));
  LUT1 #(
    .INIT(2'h1)) 
    \TX_DATA[0]_i_1 
       (.I0(TX_DATA[0]),
        .O(\TX_DATA[0]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \TX_DATA_VALID[0]_i_1 
       (.I0(TX_DATA_VALID[0]),
        .O(\TX_DATA_VALID[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \TX_DATA_VALID[1]_i_1 
       (.I0(TX_DATA_VALID[0]),
        .I1(TX_DATA_VALID[1]),
        .O(\TX_DATA_VALID[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \TX_DATA_VALID[2]_i_1 
       (.I0(TX_DATA_VALID[0]),
        .I1(TX_DATA_VALID[1]),
        .I2(TX_DATA_VALID[2]),
        .O(\TX_DATA_VALID[2]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h7F80)) 
    \TX_DATA_VALID[3]_i_1 
       (.I0(TX_DATA_VALID[1]),
        .I1(TX_DATA_VALID[0]),
        .I2(TX_DATA_VALID[2]),
        .I3(TX_DATA_VALID[3]),
        .O(\TX_DATA_VALID[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \TX_DATA_VALID[4]_i_1 
       (.I0(TX_DATA_VALID[2]),
        .I1(TX_DATA_VALID[0]),
        .I2(TX_DATA_VALID[1]),
        .I3(TX_DATA_VALID[3]),
        .I4(TX_DATA_VALID[4]),
        .O(\TX_DATA_VALID[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \TX_DATA_VALID[5]_i_1 
       (.I0(TX_DATA_VALID[3]),
        .I1(TX_DATA_VALID[1]),
        .I2(TX_DATA_VALID[0]),
        .I3(TX_DATA_VALID[2]),
        .I4(TX_DATA_VALID[4]),
        .I5(TX_DATA_VALID[5]),
        .O(\TX_DATA_VALID[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \TX_DATA_VALID[6]_i_1 
       (.I0(\TX_DATA_VALID[7]_i_2_n_0 ),
        .I1(TX_DATA_VALID[6]),
        .O(\TX_DATA_VALID[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \TX_DATA_VALID[7]_i_1 
       (.I0(\TX_DATA_VALID[7]_i_2_n_0 ),
        .I1(TX_DATA_VALID[6]),
        .I2(TX_DATA_VALID[7]),
        .O(\TX_DATA_VALID[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \TX_DATA_VALID[7]_i_2 
       (.I0(TX_DATA_VALID[5]),
        .I1(TX_DATA_VALID[3]),
        .I2(TX_DATA_VALID[1]),
        .I3(TX_DATA_VALID[0]),
        .I4(TX_DATA_VALID[2]),
        .I5(TX_DATA_VALID[4]),
        .O(\TX_DATA_VALID[7]_i_2_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[0]_i_1_n_0 ),
        .Q(TX_DATA_VALID[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[1]_i_1_n_0 ),
        .Q(TX_DATA_VALID[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[2]_i_1_n_0 ),
        .Q(TX_DATA_VALID[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[3]_i_1_n_0 ),
        .Q(TX_DATA_VALID[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[4]_i_1_n_0 ),
        .Q(TX_DATA_VALID[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[5]_i_1_n_0 ),
        .Q(TX_DATA_VALID[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[6]_i_1_n_0 ),
        .Q(TX_DATA_VALID[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_VALID[7]_i_1_n_0 ),
        .Q(TX_DATA_VALID[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA[0]_i_1_n_0 ),
        .Q(TX_DATA[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_14 ),
        .Q(TX_DATA[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[11] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_13 ),
        .Q(TX_DATA[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[12] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_12 ),
        .Q(TX_DATA[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[13] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_11 ),
        .Q(TX_DATA[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[14] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_10 ),
        .Q(TX_DATA[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[15] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_9 ),
        .Q(TX_DATA[15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[16] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_8 ),
        .Q(TX_DATA[16]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[16]_i_1 
       (.CI(\TX_DATA_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[16]_i_1_n_0 ,\TX_DATA_reg[16]_i_1_n_1 ,\TX_DATA_reg[16]_i_1_n_2 ,\TX_DATA_reg[16]_i_1_n_3 ,\TX_DATA_reg[16]_i_1_n_4 ,\TX_DATA_reg[16]_i_1_n_5 ,\TX_DATA_reg[16]_i_1_n_6 ,\TX_DATA_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[16]_i_1_n_8 ,\TX_DATA_reg[16]_i_1_n_9 ,\TX_DATA_reg[16]_i_1_n_10 ,\TX_DATA_reg[16]_i_1_n_11 ,\TX_DATA_reg[16]_i_1_n_12 ,\TX_DATA_reg[16]_i_1_n_13 ,\TX_DATA_reg[16]_i_1_n_14 ,\TX_DATA_reg[16]_i_1_n_15 }),
        .S(TX_DATA[16:9]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[17] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_15 ),
        .Q(TX_DATA[17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[18] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_14 ),
        .Q(TX_DATA[18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[19] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_13 ),
        .Q(TX_DATA[19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_15 ),
        .Q(TX_DATA[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[20] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_12 ),
        .Q(TX_DATA[20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[21] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_11 ),
        .Q(TX_DATA[21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[22] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_10 ),
        .Q(TX_DATA[22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[23] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_9 ),
        .Q(TX_DATA[23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[24] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[24]_i_1_n_8 ),
        .Q(TX_DATA[24]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[24]_i_1 
       (.CI(\TX_DATA_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[24]_i_1_n_0 ,\TX_DATA_reg[24]_i_1_n_1 ,\TX_DATA_reg[24]_i_1_n_2 ,\TX_DATA_reg[24]_i_1_n_3 ,\TX_DATA_reg[24]_i_1_n_4 ,\TX_DATA_reg[24]_i_1_n_5 ,\TX_DATA_reg[24]_i_1_n_6 ,\TX_DATA_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[24]_i_1_n_8 ,\TX_DATA_reg[24]_i_1_n_9 ,\TX_DATA_reg[24]_i_1_n_10 ,\TX_DATA_reg[24]_i_1_n_11 ,\TX_DATA_reg[24]_i_1_n_12 ,\TX_DATA_reg[24]_i_1_n_13 ,\TX_DATA_reg[24]_i_1_n_14 ,\TX_DATA_reg[24]_i_1_n_15 }),
        .S(TX_DATA[24:17]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[25] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_15 ),
        .Q(TX_DATA[25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[26] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_14 ),
        .Q(TX_DATA[26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[27] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_13 ),
        .Q(TX_DATA[27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[28] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_12 ),
        .Q(TX_DATA[28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[29] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_11 ),
        .Q(TX_DATA[29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_14 ),
        .Q(TX_DATA[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[30] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_10 ),
        .Q(TX_DATA[30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[31] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_9 ),
        .Q(TX_DATA[31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[32] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[32]_i_1_n_8 ),
        .Q(TX_DATA[32]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[32]_i_1 
       (.CI(\TX_DATA_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[32]_i_1_n_0 ,\TX_DATA_reg[32]_i_1_n_1 ,\TX_DATA_reg[32]_i_1_n_2 ,\TX_DATA_reg[32]_i_1_n_3 ,\TX_DATA_reg[32]_i_1_n_4 ,\TX_DATA_reg[32]_i_1_n_5 ,\TX_DATA_reg[32]_i_1_n_6 ,\TX_DATA_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[32]_i_1_n_8 ,\TX_DATA_reg[32]_i_1_n_9 ,\TX_DATA_reg[32]_i_1_n_10 ,\TX_DATA_reg[32]_i_1_n_11 ,\TX_DATA_reg[32]_i_1_n_12 ,\TX_DATA_reg[32]_i_1_n_13 ,\TX_DATA_reg[32]_i_1_n_14 ,\TX_DATA_reg[32]_i_1_n_15 }),
        .S(TX_DATA[32:25]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[33] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_15 ),
        .Q(TX_DATA[33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[34] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_14 ),
        .Q(TX_DATA[34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[35] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_13 ),
        .Q(TX_DATA[35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[36] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_12 ),
        .Q(TX_DATA[36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[37] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_11 ),
        .Q(TX_DATA[37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[38] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_10 ),
        .Q(TX_DATA[38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[39] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_9 ),
        .Q(TX_DATA[39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_13 ),
        .Q(TX_DATA[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[40] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[40]_i_1_n_8 ),
        .Q(TX_DATA[40]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[40]_i_1 
       (.CI(\TX_DATA_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[40]_i_1_n_0 ,\TX_DATA_reg[40]_i_1_n_1 ,\TX_DATA_reg[40]_i_1_n_2 ,\TX_DATA_reg[40]_i_1_n_3 ,\TX_DATA_reg[40]_i_1_n_4 ,\TX_DATA_reg[40]_i_1_n_5 ,\TX_DATA_reg[40]_i_1_n_6 ,\TX_DATA_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[40]_i_1_n_8 ,\TX_DATA_reg[40]_i_1_n_9 ,\TX_DATA_reg[40]_i_1_n_10 ,\TX_DATA_reg[40]_i_1_n_11 ,\TX_DATA_reg[40]_i_1_n_12 ,\TX_DATA_reg[40]_i_1_n_13 ,\TX_DATA_reg[40]_i_1_n_14 ,\TX_DATA_reg[40]_i_1_n_15 }),
        .S(TX_DATA[40:33]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[41] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_15 ),
        .Q(TX_DATA[41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[42] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_14 ),
        .Q(TX_DATA[42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[43] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_13 ),
        .Q(TX_DATA[43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[44] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_12 ),
        .Q(TX_DATA[44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[45] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_11 ),
        .Q(TX_DATA[45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[46] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_10 ),
        .Q(TX_DATA[46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[47] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_9 ),
        .Q(TX_DATA[47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[48] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[48]_i_1_n_8 ),
        .Q(TX_DATA[48]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[48]_i_1 
       (.CI(\TX_DATA_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[48]_i_1_n_0 ,\TX_DATA_reg[48]_i_1_n_1 ,\TX_DATA_reg[48]_i_1_n_2 ,\TX_DATA_reg[48]_i_1_n_3 ,\TX_DATA_reg[48]_i_1_n_4 ,\TX_DATA_reg[48]_i_1_n_5 ,\TX_DATA_reg[48]_i_1_n_6 ,\TX_DATA_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[48]_i_1_n_8 ,\TX_DATA_reg[48]_i_1_n_9 ,\TX_DATA_reg[48]_i_1_n_10 ,\TX_DATA_reg[48]_i_1_n_11 ,\TX_DATA_reg[48]_i_1_n_12 ,\TX_DATA_reg[48]_i_1_n_13 ,\TX_DATA_reg[48]_i_1_n_14 ,\TX_DATA_reg[48]_i_1_n_15 }),
        .S(TX_DATA[48:41]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[49] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_15 ),
        .Q(TX_DATA[49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_12 ),
        .Q(TX_DATA[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[50] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_14 ),
        .Q(TX_DATA[50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[51] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_13 ),
        .Q(TX_DATA[51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[52] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_12 ),
        .Q(TX_DATA[52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[53] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_11 ),
        .Q(TX_DATA[53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[54] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_10 ),
        .Q(TX_DATA[54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[55] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_9 ),
        .Q(TX_DATA[55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[56] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[56]_i_1_n_8 ),
        .Q(TX_DATA[56]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[56]_i_1 
       (.CI(\TX_DATA_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[56]_i_1_n_0 ,\TX_DATA_reg[56]_i_1_n_1 ,\TX_DATA_reg[56]_i_1_n_2 ,\TX_DATA_reg[56]_i_1_n_3 ,\TX_DATA_reg[56]_i_1_n_4 ,\TX_DATA_reg[56]_i_1_n_5 ,\TX_DATA_reg[56]_i_1_n_6 ,\TX_DATA_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[56]_i_1_n_8 ,\TX_DATA_reg[56]_i_1_n_9 ,\TX_DATA_reg[56]_i_1_n_10 ,\TX_DATA_reg[56]_i_1_n_11 ,\TX_DATA_reg[56]_i_1_n_12 ,\TX_DATA_reg[56]_i_1_n_13 ,\TX_DATA_reg[56]_i_1_n_14 ,\TX_DATA_reg[56]_i_1_n_15 }),
        .S(TX_DATA[56:49]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[57] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_15 ),
        .Q(TX_DATA[57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[58] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_14 ),
        .Q(TX_DATA[58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[59] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_13 ),
        .Q(TX_DATA[59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_11 ),
        .Q(TX_DATA[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[60] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_12 ),
        .Q(TX_DATA[60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[61] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_11 ),
        .Q(TX_DATA[61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[62] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_10 ),
        .Q(TX_DATA[62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[63] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[63]_i_1_n_9 ),
        .Q(TX_DATA[63]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[63]_i_1 
       (.CI(\TX_DATA_reg[56]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_TX_DATA_reg[63]_i_1_CO_UNCONNECTED [7:6],\TX_DATA_reg[63]_i_1_n_2 ,\TX_DATA_reg[63]_i_1_n_3 ,\TX_DATA_reg[63]_i_1_n_4 ,\TX_DATA_reg[63]_i_1_n_5 ,\TX_DATA_reg[63]_i_1_n_6 ,\TX_DATA_reg[63]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_TX_DATA_reg[63]_i_1_O_UNCONNECTED [7],\TX_DATA_reg[63]_i_1_n_9 ,\TX_DATA_reg[63]_i_1_n_10 ,\TX_DATA_reg[63]_i_1_n_11 ,\TX_DATA_reg[63]_i_1_n_12 ,\TX_DATA_reg[63]_i_1_n_13 ,\TX_DATA_reg[63]_i_1_n_14 ,\TX_DATA_reg[63]_i_1_n_15 }),
        .S({1'b0,TX_DATA[63:57]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_10 ),
        .Q(TX_DATA[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_9 ),
        .Q(TX_DATA[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[8]_i_1_n_8 ),
        .Q(TX_DATA[8]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \TX_DATA_reg[8]_i_1 
       (.CI(TX_DATA[0]),
        .CI_TOP(1'b0),
        .CO({\TX_DATA_reg[8]_i_1_n_0 ,\TX_DATA_reg[8]_i_1_n_1 ,\TX_DATA_reg[8]_i_1_n_2 ,\TX_DATA_reg[8]_i_1_n_3 ,\TX_DATA_reg[8]_i_1_n_4 ,\TX_DATA_reg[8]_i_1_n_5 ,\TX_DATA_reg[8]_i_1_n_6 ,\TX_DATA_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\TX_DATA_reg[8]_i_1_n_8 ,\TX_DATA_reg[8]_i_1_n_9 ,\TX_DATA_reg[8]_i_1_n_10 ,\TX_DATA_reg[8]_i_1_n_11 ,\TX_DATA_reg[8]_i_1_n_12 ,\TX_DATA_reg[8]_i_1_n_13 ,\TX_DATA_reg[8]_i_1_n_14 ,\TX_DATA_reg[8]_i_1_n_15 }),
        .S(TX_DATA[8:1]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_DATA_reg[16]_i_1_n_15 ),
        .Q(TX_DATA[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h1)) 
    \TX_IFG_DELAY[0]_i_1 
       (.I0(TX_IFG_DELAY[0]),
        .O(\TX_IFG_DELAY[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \TX_IFG_DELAY[1]_i_1 
       (.I0(TX_IFG_DELAY[0]),
        .I1(TX_IFG_DELAY[1]),
        .O(\TX_IFG_DELAY[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \TX_IFG_DELAY[2]_i_1 
       (.I0(TX_IFG_DELAY[0]),
        .I1(TX_IFG_DELAY[1]),
        .I2(TX_IFG_DELAY[2]),
        .O(\TX_IFG_DELAY[2]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h7F80)) 
    \TX_IFG_DELAY[3]_i_1 
       (.I0(TX_IFG_DELAY[1]),
        .I1(TX_IFG_DELAY[0]),
        .I2(TX_IFG_DELAY[2]),
        .I3(TX_IFG_DELAY[3]),
        .O(\TX_IFG_DELAY[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \TX_IFG_DELAY[4]_i_1 
       (.I0(TX_IFG_DELAY[2]),
        .I1(TX_IFG_DELAY[0]),
        .I2(TX_IFG_DELAY[1]),
        .I3(TX_IFG_DELAY[3]),
        .I4(TX_IFG_DELAY[4]),
        .O(\TX_IFG_DELAY[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \TX_IFG_DELAY[5]_i_1 
       (.I0(TX_IFG_DELAY[3]),
        .I1(TX_IFG_DELAY[1]),
        .I2(TX_IFG_DELAY[0]),
        .I3(TX_IFG_DELAY[2]),
        .I4(TX_IFG_DELAY[4]),
        .I5(TX_IFG_DELAY[5]),
        .O(\TX_IFG_DELAY[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \TX_IFG_DELAY[6]_i_1 
       (.I0(\TX_IFG_DELAY[7]_i_2_n_0 ),
        .I1(TX_IFG_DELAY[6]),
        .O(\TX_IFG_DELAY[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \TX_IFG_DELAY[7]_i_1 
       (.I0(\TX_IFG_DELAY[7]_i_2_n_0 ),
        .I1(TX_IFG_DELAY[6]),
        .I2(TX_IFG_DELAY[7]),
        .O(\TX_IFG_DELAY[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \TX_IFG_DELAY[7]_i_2 
       (.I0(TX_IFG_DELAY[5]),
        .I1(TX_IFG_DELAY[3]),
        .I2(TX_IFG_DELAY[1]),
        .I3(TX_IFG_DELAY[0]),
        .I4(TX_IFG_DELAY[2]),
        .I5(TX_IFG_DELAY[4]),
        .O(\TX_IFG_DELAY[7]_i_2_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[0]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[1]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[2]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[3]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[4]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[5]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[6]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \TX_IFG_DELAY_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\TX_IFG_DELAY[7]_i_1_n_0 ),
        .Q(TX_IFG_DELAY[7]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h2)) 
    TX_START_inst
       (.I0(wdata[6]),
        .O(TX_START));
  LUT1 #(
    .INIT(2'h2)) 
    TX_UNDERRUN_inst
       (.I0(dat_i),
        .O(TX_UNDERRUN));
  switch_elements_cfg_crc \activity_blocks[0].dutA 
       (.Q(dat_o_vec),
        .clk_i(rxclk_out),
        .\dat_o_reg[0]_0 (dat_i),
        .out(crc_en),
        .rst_i(rst_i));
  switch_elements_simple_spi_top \activity_blocks[0].dutB 
       (.E(\activity_blocks[0].dutH_n_0 ),
        .ack_o(ack_o),
        .clk_i(rxclk_out),
        .dat_i(dat_i_vec),
        .dat_o(dat_o),
        .\dat_o_reg[3]_0 (adr_i),
        .in0(inta_o),
        .out(we_i),
        .rst_i(rst_i),
        .sck_o(sck_o),
        .\sper_reg[0]_0 (cyc_i),
        .\sper_reg[0]_1 (stb_i),
        .treg(mosi_o),
        .\treg_reg[0]_0 (miso_i));
  switch_elements_management_top \activity_blocks[0].dutC 
       (.CLK(mdc),
        .cfgRxRegData(cfgRxRegData),
        .cfgTxRegData(cfgTxRegData),
        .clk_i(rxclk_out),
        .in0(mgmt_miim_rdy),
        .mdio_i(mdio),
        .mgmt_rd_data(mgmt_rd_data),
        .mgmt_wr_data(mgmt_wr_data),
        .out(mgmt_addr),
        .\recv_config0_reg[0] (mgmt_opcode[1]),
        .rst_i(rst_i),
        .rxStatRegPlus({rxStatRegPlus[18:7],dat_i_vec[6:0]}),
        .\stat_rd_data_reg[63] (mgmt_req),
        .\stat_rd_data_reg[63]_0 (mgmt_miim_sel),
        .txStatRegPlus(txStatRegPlus[14:0]));
  switch_elements_rxReceiveEngine \activity_blocks[0].dutD 
       (.D(xgmii_rxd),
        .Q(rxTxLinkFault_vec),
        .\cfgRxRegData_reg[52]_0 (cfgRxRegData_in[52:48]),
        .clk_i(rxclk_out),
        .in0({rxStatRegPlus[17:14],rxStatRegPlus[11],rxStatRegPlus[8:0]}),
        .rst_i(rst_i),
        .rxCfgofRS(rxCfgofRS),
        .rx_bad_frame(rx_bad_frame),
        .rx_data(rx_data),
        .rx_data_valid(rx_data_valid),
        .rx_good_frame(rx_good_frame),
        .\rxc4_in_tmp_reg[3] (xgmii_rxc),
        .rxclk_180(rxclk_180));
  switch_elements_manchesterWireless \activity_blocks[0].dutE 
       (.clk_i(rxclk_out),
        .in0(recieved_debug),
        .out(data_i),
        .q_o(q_o),
        .ready_o(ready_o),
        .rst_i(rst_i),
        .waitforstart_rdy(waitforstart_rdy));
  switch_elements_LPF3x8 \activity_blocks[0].dutG 
       (.DI(DI),
        .DO(DO),
        .E(\activity_blocks[0].dutH_n_0 ),
        .FREQ(FREQ),
        .clk_i(rxclk_out),
        .d4_30(d4_30),
        .\d4_4_reg[15]_0 (activity_blocks_c_11_n_0),
        .out(EF),
        .rst_i(rst_i));
  switch_elements_TRANSMIT_TOP \activity_blocks[0].dutH 
       (.\DELAY_ACK_reg[7]_0 (TX_IFG_DELAY),
        .E(\activity_blocks[0].dutH_n_0 ),
        .FC_TRANS_PAUSEDATA(FC_TRANS_PAUSEDATA),
        .FC_TRANS_PAUSEVAL(FC_TRANS_PAUSEVAL),
        .I94(FC_TX_PAUSEDATA),
        .TXC(TXC),
        .TXD(TXD),
        .TXSTATREGPLUS(txStatRegPlus),
        .TX_ACK(TX_ACK),
        .TX_CFG_REG_VALID(TX_CFG_REG_VALID),
        .TX_CFG_REG_VALUE({TX_CFG_REG_VALUE[31],TX_CFG_REG_VALUE[29],TX_CFG_REG_VALUE[27],TX_CFG_REG_VALUE[25]}),
        .TX_DATA(TX_DATA),
        .\TX_DATA_VALID_REG_reg[7]_0 (TX_DATA_VALID),
        .TX_STATS_VALID(TX_STATS_VALID),
        .apply_pause_delay_reg_0(FC_TX_PAUSEVALID),
        .clk_i(rxclk_out),
        .load_final_CRC_reg_0(activity_blocks_c_8_n_0),
        .out(TX_START),
        .rst_i(rst_i),
        .tx_undderrun_int_reg_0(TX_UNDERRUN));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(1'b1),
        .Q(activity_blocks_c_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_0
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_n_0),
        .Q(activity_blocks_c_0_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_1
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_0_n_0),
        .Q(activity_blocks_c_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_10
       (.C(rxclk_out),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_c_9_n_0),
        .Q(activity_blocks_c_10_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_11
       (.C(rxclk_out),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_c_10_n_0),
        .Q(activity_blocks_c_11_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_2
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_1_n_0),
        .Q(activity_blocks_c_2_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_3
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_2_n_0),
        .Q(activity_blocks_c_3_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_4
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_3_n_0),
        .Q(activity_blocks_c_4_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_5
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_4_n_0),
        .Q(activity_blocks_c_5_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_6
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_5_n_0),
        .Q(activity_blocks_c_6_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_7
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_6_n_0),
        .Q(activity_blocks_c_7_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_8
       (.C(rxclk_out),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_c_7_n_0),
        .Q(activity_blocks_c_8_n_0));
  FDCE #(
    .INIT(1'b0)) 
    activity_blocks_c_9
       (.C(rxclk_out),
        .CE(d4_30),
        .CLR(rst_i),
        .D(1'b1),
        .Q(activity_blocks_c_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    \addr[0]_i_1 
       (.I0(addr[0]),
        .O(\addr[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \addr[10]_i_1 
       (.I0(addr[8]),
        .I1(addr[6]),
        .I2(\addr[10]_i_2_n_0 ),
        .I3(addr[7]),
        .I4(addr[9]),
        .I5(addr[10]),
        .O(\addr[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \addr[10]_i_2 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[1]),
        .I3(addr[0]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\addr[10]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \addr[1]_i_1 
       (.I0(addr[0]),
        .I1(addr[1]),
        .O(\addr[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \addr[2]_i_1 
       (.I0(addr[0]),
        .I1(addr[1]),
        .I2(addr[2]),
        .O(\addr[2]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h7F80)) 
    \addr[3]_i_1 
       (.I0(addr[1]),
        .I1(addr[0]),
        .I2(addr[2]),
        .I3(addr[3]),
        .O(\addr[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \addr[4]_i_1 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .O(\addr[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \addr[5]_i_1 
       (.I0(addr[3]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[2]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\addr[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \addr[6]_i_1 
       (.I0(\addr[10]_i_2_n_0 ),
        .I1(addr[6]),
        .O(\addr[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \addr[7]_i_1 
       (.I0(\addr[10]_i_2_n_0 ),
        .I1(addr[6]),
        .I2(addr[7]),
        .O(\addr[7]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h7F80)) 
    \addr[8]_i_1 
       (.I0(addr[6]),
        .I1(\addr[10]_i_2_n_0 ),
        .I2(addr[7]),
        .I3(addr[8]),
        .O(\addr[8]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \addr[9]_i_1 
       (.I0(addr[7]),
        .I1(\addr[10]_i_2_n_0 ),
        .I2(addr[6]),
        .I3(addr[8]),
        .I4(addr[9]),
        .O(\addr[9]_i_1_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[0]_i_1_n_0 ),
        .Q(addr[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[10]_i_1_n_0 ),
        .Q(addr[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[1]_i_1_n_0 ),
        .Q(addr[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[2]_i_1_n_0 ),
        .Q(addr[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[3]_i_1_n_0 ),
        .Q(addr[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[4]_i_1_n_0 ),
        .Q(addr[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[5]_i_1_n_0 ),
        .Q(addr[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[6]_i_1_n_0 ),
        .Q(addr[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[7]_i_1_n_0 ),
        .Q(addr[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[8]_i_1_n_0 ),
        .Q(addr[8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \addr_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\addr[9]_i_1_n_0 ),
        .Q(addr[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h2)) 
    adr_i_inst
       (.I0(wdata[5]),
        .O(adr_i[1]));
  LUT1 #(
    .INIT(2'h2)) 
    adr_i_inst__0
       (.I0(wdata[4]),
        .O(adr_i[0]));
  LUT1 #(
    .INIT(2'h1)) 
    \cfgRxRegData_in[0]_i_1 
       (.I0(cfgRxRegData_in[0]),
        .O(\cfgRxRegData_in[0]_i_1_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in[0]_i_1_n_0 ),
        .Q(cfgRxRegData_in[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_14 ),
        .Q(cfgRxRegData_in[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[11] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_13 ),
        .Q(cfgRxRegData_in[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[12] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_12 ),
        .Q(cfgRxRegData_in[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[13] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_11 ),
        .Q(cfgRxRegData_in[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[14] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_10 ),
        .Q(cfgRxRegData_in[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[15] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_9 ),
        .Q(cfgRxRegData_in[15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[16] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_8 ),
        .Q(cfgRxRegData_in[16]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[16]_i_1 
       (.CI(\cfgRxRegData_in_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[16]_i_1_n_0 ,\cfgRxRegData_in_reg[16]_i_1_n_1 ,\cfgRxRegData_in_reg[16]_i_1_n_2 ,\cfgRxRegData_in_reg[16]_i_1_n_3 ,\cfgRxRegData_in_reg[16]_i_1_n_4 ,\cfgRxRegData_in_reg[16]_i_1_n_5 ,\cfgRxRegData_in_reg[16]_i_1_n_6 ,\cfgRxRegData_in_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[16]_i_1_n_8 ,\cfgRxRegData_in_reg[16]_i_1_n_9 ,\cfgRxRegData_in_reg[16]_i_1_n_10 ,\cfgRxRegData_in_reg[16]_i_1_n_11 ,\cfgRxRegData_in_reg[16]_i_1_n_12 ,\cfgRxRegData_in_reg[16]_i_1_n_13 ,\cfgRxRegData_in_reg[16]_i_1_n_14 ,\cfgRxRegData_in_reg[16]_i_1_n_15 }),
        .S(cfgRxRegData_in[16:9]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[17] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_15 ),
        .Q(cfgRxRegData_in[17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[18] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_14 ),
        .Q(cfgRxRegData_in[18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[19] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_13 ),
        .Q(cfgRxRegData_in[19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_15 ),
        .Q(cfgRxRegData_in[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[20] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_12 ),
        .Q(cfgRxRegData_in[20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[21] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_11 ),
        .Q(cfgRxRegData_in[21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[22] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_10 ),
        .Q(cfgRxRegData_in[22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[23] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_9 ),
        .Q(cfgRxRegData_in[23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[24] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[24]_i_1_n_8 ),
        .Q(cfgRxRegData_in[24]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[24]_i_1 
       (.CI(\cfgRxRegData_in_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[24]_i_1_n_0 ,\cfgRxRegData_in_reg[24]_i_1_n_1 ,\cfgRxRegData_in_reg[24]_i_1_n_2 ,\cfgRxRegData_in_reg[24]_i_1_n_3 ,\cfgRxRegData_in_reg[24]_i_1_n_4 ,\cfgRxRegData_in_reg[24]_i_1_n_5 ,\cfgRxRegData_in_reg[24]_i_1_n_6 ,\cfgRxRegData_in_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[24]_i_1_n_8 ,\cfgRxRegData_in_reg[24]_i_1_n_9 ,\cfgRxRegData_in_reg[24]_i_1_n_10 ,\cfgRxRegData_in_reg[24]_i_1_n_11 ,\cfgRxRegData_in_reg[24]_i_1_n_12 ,\cfgRxRegData_in_reg[24]_i_1_n_13 ,\cfgRxRegData_in_reg[24]_i_1_n_14 ,\cfgRxRegData_in_reg[24]_i_1_n_15 }),
        .S(cfgRxRegData_in[24:17]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[25] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_15 ),
        .Q(cfgRxRegData_in[25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[26] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_14 ),
        .Q(cfgRxRegData_in[26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[27] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_13 ),
        .Q(cfgRxRegData_in[27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[28] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_12 ),
        .Q(cfgRxRegData_in[28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[29] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_11 ),
        .Q(cfgRxRegData_in[29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_14 ),
        .Q(cfgRxRegData_in[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[30] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_10 ),
        .Q(cfgRxRegData_in[30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[31] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_9 ),
        .Q(cfgRxRegData_in[31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[32] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[32]_i_1_n_8 ),
        .Q(cfgRxRegData_in[32]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[32]_i_1 
       (.CI(\cfgRxRegData_in_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[32]_i_1_n_0 ,\cfgRxRegData_in_reg[32]_i_1_n_1 ,\cfgRxRegData_in_reg[32]_i_1_n_2 ,\cfgRxRegData_in_reg[32]_i_1_n_3 ,\cfgRxRegData_in_reg[32]_i_1_n_4 ,\cfgRxRegData_in_reg[32]_i_1_n_5 ,\cfgRxRegData_in_reg[32]_i_1_n_6 ,\cfgRxRegData_in_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[32]_i_1_n_8 ,\cfgRxRegData_in_reg[32]_i_1_n_9 ,\cfgRxRegData_in_reg[32]_i_1_n_10 ,\cfgRxRegData_in_reg[32]_i_1_n_11 ,\cfgRxRegData_in_reg[32]_i_1_n_12 ,\cfgRxRegData_in_reg[32]_i_1_n_13 ,\cfgRxRegData_in_reg[32]_i_1_n_14 ,\cfgRxRegData_in_reg[32]_i_1_n_15 }),
        .S(cfgRxRegData_in[32:25]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[33] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_15 ),
        .Q(cfgRxRegData_in[33]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[34] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_14 ),
        .Q(cfgRxRegData_in[34]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[35] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_13 ),
        .Q(cfgRxRegData_in[35]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[36] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_12 ),
        .Q(cfgRxRegData_in[36]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[37] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_11 ),
        .Q(cfgRxRegData_in[37]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[38] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_10 ),
        .Q(cfgRxRegData_in[38]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[39] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_9 ),
        .Q(cfgRxRegData_in[39]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_13 ),
        .Q(cfgRxRegData_in[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[40] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[40]_i_1_n_8 ),
        .Q(cfgRxRegData_in[40]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[40]_i_1 
       (.CI(\cfgRxRegData_in_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[40]_i_1_n_0 ,\cfgRxRegData_in_reg[40]_i_1_n_1 ,\cfgRxRegData_in_reg[40]_i_1_n_2 ,\cfgRxRegData_in_reg[40]_i_1_n_3 ,\cfgRxRegData_in_reg[40]_i_1_n_4 ,\cfgRxRegData_in_reg[40]_i_1_n_5 ,\cfgRxRegData_in_reg[40]_i_1_n_6 ,\cfgRxRegData_in_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[40]_i_1_n_8 ,\cfgRxRegData_in_reg[40]_i_1_n_9 ,\cfgRxRegData_in_reg[40]_i_1_n_10 ,\cfgRxRegData_in_reg[40]_i_1_n_11 ,\cfgRxRegData_in_reg[40]_i_1_n_12 ,\cfgRxRegData_in_reg[40]_i_1_n_13 ,\cfgRxRegData_in_reg[40]_i_1_n_14 ,\cfgRxRegData_in_reg[40]_i_1_n_15 }),
        .S(cfgRxRegData_in[40:33]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[41] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_15 ),
        .Q(cfgRxRegData_in[41]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[42] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_14 ),
        .Q(cfgRxRegData_in[42]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[43] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_13 ),
        .Q(cfgRxRegData_in[43]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[44] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_12 ),
        .Q(cfgRxRegData_in[44]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[45] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_11 ),
        .Q(cfgRxRegData_in[45]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[46] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_10 ),
        .Q(cfgRxRegData_in[46]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[47] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_9 ),
        .Q(cfgRxRegData_in[47]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[48] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[48]_i_1_n_8 ),
        .Q(cfgRxRegData_in[48]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[48]_i_1 
       (.CI(\cfgRxRegData_in_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[48]_i_1_n_0 ,\cfgRxRegData_in_reg[48]_i_1_n_1 ,\cfgRxRegData_in_reg[48]_i_1_n_2 ,\cfgRxRegData_in_reg[48]_i_1_n_3 ,\cfgRxRegData_in_reg[48]_i_1_n_4 ,\cfgRxRegData_in_reg[48]_i_1_n_5 ,\cfgRxRegData_in_reg[48]_i_1_n_6 ,\cfgRxRegData_in_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[48]_i_1_n_8 ,\cfgRxRegData_in_reg[48]_i_1_n_9 ,\cfgRxRegData_in_reg[48]_i_1_n_10 ,\cfgRxRegData_in_reg[48]_i_1_n_11 ,\cfgRxRegData_in_reg[48]_i_1_n_12 ,\cfgRxRegData_in_reg[48]_i_1_n_13 ,\cfgRxRegData_in_reg[48]_i_1_n_14 ,\cfgRxRegData_in_reg[48]_i_1_n_15 }),
        .S(cfgRxRegData_in[48:41]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[49] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_15 ),
        .Q(cfgRxRegData_in[49]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_12 ),
        .Q(cfgRxRegData_in[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[50] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_14 ),
        .Q(cfgRxRegData_in[50]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[51] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_13 ),
        .Q(cfgRxRegData_in[51]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[52] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_12 ),
        .Q(cfgRxRegData_in[52]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[53] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_11 ),
        .Q(cfgRxRegData_in[53]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[54] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_10 ),
        .Q(cfgRxRegData_in[54]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[55] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_9 ),
        .Q(cfgRxRegData_in[55]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[56] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[56]_i_1_n_8 ),
        .Q(cfgRxRegData_in[56]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[56]_i_1 
       (.CI(\cfgRxRegData_in_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[56]_i_1_n_0 ,\cfgRxRegData_in_reg[56]_i_1_n_1 ,\cfgRxRegData_in_reg[56]_i_1_n_2 ,\cfgRxRegData_in_reg[56]_i_1_n_3 ,\cfgRxRegData_in_reg[56]_i_1_n_4 ,\cfgRxRegData_in_reg[56]_i_1_n_5 ,\cfgRxRegData_in_reg[56]_i_1_n_6 ,\cfgRxRegData_in_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[56]_i_1_n_8 ,\cfgRxRegData_in_reg[56]_i_1_n_9 ,\cfgRxRegData_in_reg[56]_i_1_n_10 ,\cfgRxRegData_in_reg[56]_i_1_n_11 ,\cfgRxRegData_in_reg[56]_i_1_n_12 ,\cfgRxRegData_in_reg[56]_i_1_n_13 ,\cfgRxRegData_in_reg[56]_i_1_n_14 ,\cfgRxRegData_in_reg[56]_i_1_n_15 }),
        .S(cfgRxRegData_in[56:49]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[57] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_15 ),
        .Q(cfgRxRegData_in[57]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[58] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_14 ),
        .Q(cfgRxRegData_in[58]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[59] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_13 ),
        .Q(cfgRxRegData_in[59]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_11 ),
        .Q(cfgRxRegData_in[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[60] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_12 ),
        .Q(cfgRxRegData_in[60]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[61] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_11 ),
        .Q(cfgRxRegData_in[61]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[62] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_10 ),
        .Q(cfgRxRegData_in[62]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[63] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_9 ),
        .Q(cfgRxRegData_in[63]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[64] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[64]_i_1_n_8 ),
        .Q(cfgRxRegData_in[64]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[64]_i_1 
       (.CI(\cfgRxRegData_in_reg[56]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_cfgRxRegData_in_reg[64]_i_1_CO_UNCONNECTED [7],\cfgRxRegData_in_reg[64]_i_1_n_1 ,\cfgRxRegData_in_reg[64]_i_1_n_2 ,\cfgRxRegData_in_reg[64]_i_1_n_3 ,\cfgRxRegData_in_reg[64]_i_1_n_4 ,\cfgRxRegData_in_reg[64]_i_1_n_5 ,\cfgRxRegData_in_reg[64]_i_1_n_6 ,\cfgRxRegData_in_reg[64]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[64]_i_1_n_8 ,\cfgRxRegData_in_reg[64]_i_1_n_9 ,\cfgRxRegData_in_reg[64]_i_1_n_10 ,\cfgRxRegData_in_reg[64]_i_1_n_11 ,\cfgRxRegData_in_reg[64]_i_1_n_12 ,\cfgRxRegData_in_reg[64]_i_1_n_13 ,\cfgRxRegData_in_reg[64]_i_1_n_14 ,\cfgRxRegData_in_reg[64]_i_1_n_15 }),
        .S(cfgRxRegData_in[64:57]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_10 ),
        .Q(cfgRxRegData_in[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_9 ),
        .Q(cfgRxRegData_in[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[8]_i_1_n_8 ),
        .Q(cfgRxRegData_in[8]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \cfgRxRegData_in_reg[8]_i_1 
       (.CI(cfgRxRegData_in[0]),
        .CI_TOP(1'b0),
        .CO({\cfgRxRegData_in_reg[8]_i_1_n_0 ,\cfgRxRegData_in_reg[8]_i_1_n_1 ,\cfgRxRegData_in_reg[8]_i_1_n_2 ,\cfgRxRegData_in_reg[8]_i_1_n_3 ,\cfgRxRegData_in_reg[8]_i_1_n_4 ,\cfgRxRegData_in_reg[8]_i_1_n_5 ,\cfgRxRegData_in_reg[8]_i_1_n_6 ,\cfgRxRegData_in_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\cfgRxRegData_in_reg[8]_i_1_n_8 ,\cfgRxRegData_in_reg[8]_i_1_n_9 ,\cfgRxRegData_in_reg[8]_i_1_n_10 ,\cfgRxRegData_in_reg[8]_i_1_n_11 ,\cfgRxRegData_in_reg[8]_i_1_n_12 ,\cfgRxRegData_in_reg[8]_i_1_n_13 ,\cfgRxRegData_in_reg[8]_i_1_n_14 ,\cfgRxRegData_in_reg[8]_i_1_n_15 }),
        .S(cfgRxRegData_in[8:1]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \cfgRxRegData_in_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\cfgRxRegData_in_reg[16]_i_1_n_15 ),
        .Q(cfgRxRegData_in[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h2)) 
    cyc_i_inst
       (.I0(wdata[2]),
        .O(cyc_i));
  LUT1 #(
    .INIT(2'h2)) 
    dat_i_vec_inst
       (.I0(wdata[1]),
        .O(dat_i_vec[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(outputs[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(outputs[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(rdata[13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(rdata[12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(rdata[11]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(rdata[10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(rdata[9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(rdata[8]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(rdata[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(rdata[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(rdata[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(rdata[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(outputs[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(rdata[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(rdata[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(rdata[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(rdata[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(rxStatRegPlus[18]));
  LUT1 #(
    .INIT(2'h2)) 
    i_25
       (.I0(1'b0),
        .O(rxStatRegPlus[13]));
  LUT1 #(
    .INIT(2'h2)) 
    i_26
       (.I0(1'b0),
        .O(rxStatRegPlus[12]));
  LUT1 #(
    .INIT(2'h2)) 
    i_27
       (.I0(1'b0),
        .O(rxStatRegPlus[10]));
  LUT1 #(
    .INIT(2'h2)) 
    i_28
       (.I0(1'b0),
        .O(rxStatRegPlus[9]));
  LUT1 #(
    .INIT(2'h2)) 
    i_29
       (.I0(1'b0),
        .O(data_i));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(outputs[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_30
       (.I0(1'b0),
        .O(mdio));
  LUT1 #(
    .INIT(2'h2)) 
    i_31
       (.I0(1'b0),
        .O(run_out));
  LUT1 #(
    .INIT(2'h2)) 
    i_32
       (.I0(1'b0),
        .O(rst_syn));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(outputs[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(outputs[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(outputs[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(outputs[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(rdata[15]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(rdata[14]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \info_o[0]_INST_0 
       (.I0(outputs[0]),
        .I1(rdata[0]),
        .I2(mosi_o),
        .I3(q_o[0]),
        .I4(\info_o[0]_INST_0_i_1_n_0 ),
        .O(info_o[0]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[0]_INST_0_i_1 
       (.I0(rx_data[0]),
        .I1(DO[0]),
        .I2(dat_o[0]),
        .I3(TXD[0]),
        .O(\info_o[0]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[10]_INST_0 
       (.I0(rx_data[10]),
        .I1(DO[10]),
        .I2(rdata[10]),
        .I3(TXD[10]),
        .O(info_o[10]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[11]_INST_0 
       (.I0(rx_data[11]),
        .I1(DO[11]),
        .I2(rdata[11]),
        .I3(TXD[11]),
        .O(info_o[11]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[12]_INST_0 
       (.I0(rx_data[12]),
        .I1(DO[12]),
        .I2(rdata[12]),
        .I3(TXD[12]),
        .O(info_o[12]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[13]_INST_0 
       (.I0(rx_data[13]),
        .I1(DO[13]),
        .I2(rdata[13]),
        .I3(TXD[13]),
        .O(info_o[13]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[14]_INST_0 
       (.I0(rx_data[14]),
        .I1(DO[14]),
        .I2(rdata[14]),
        .I3(TXD[14]),
        .O(info_o[14]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[15]_INST_0 
       (.I0(rx_data[15]),
        .I1(DO[15]),
        .I2(rdata[15]),
        .I3(TXD[15]),
        .O(info_o[15]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[16]_INST_0 
       (.I0(rx_data[16]),
        .I1(TXD[16]),
        .I2(cfgRxRegData[16]),
        .O(info_o[16]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[17]_INST_0 
       (.I0(rx_data[17]),
        .I1(TXD[17]),
        .I2(cfgRxRegData[17]),
        .O(info_o[17]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[18]_INST_0 
       (.I0(rx_data[18]),
        .I1(TXD[18]),
        .I2(cfgRxRegData[18]),
        .O(info_o[18]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[19]_INST_0 
       (.I0(rx_data[19]),
        .I1(TXD[19]),
        .I2(cfgRxRegData[19]),
        .O(info_o[19]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[1]_INST_0 
       (.I0(rdata[1]),
        .I1(outputs[1]),
        .I2(TXD[1]),
        .I3(dat_o[1]),
        .I4(DO[1]),
        .I5(rx_data[1]),
        .O(info_o[1]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[20]_INST_0 
       (.I0(rx_data[20]),
        .I1(TXD[20]),
        .I2(cfgRxRegData[20]),
        .O(info_o[20]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[21]_INST_0 
       (.I0(rx_data[21]),
        .I1(TXD[21]),
        .I2(cfgRxRegData[21]),
        .O(info_o[21]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[22]_INST_0 
       (.I0(rx_data[22]),
        .I1(TXD[22]),
        .I2(cfgRxRegData[22]),
        .O(info_o[22]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[23]_INST_0 
       (.I0(rx_data[23]),
        .I1(TXD[23]),
        .I2(cfgRxRegData[23]),
        .O(info_o[23]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[24]_INST_0 
       (.I0(rx_data[24]),
        .I1(TXD[24]),
        .I2(cfgRxRegData[24]),
        .O(info_o[24]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[25]_INST_0 
       (.I0(rx_data[25]),
        .I1(TXD[25]),
        .I2(cfgRxRegData[25]),
        .O(info_o[25]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[26]_INST_0 
       (.I0(rx_data[26]),
        .I1(TXD[26]),
        .I2(cfgRxRegData[26]),
        .O(info_o[26]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[27]_INST_0 
       (.I0(rx_data[27]),
        .I1(TXD[27]),
        .I2(cfgRxRegData[27]),
        .O(info_o[27]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[28]_INST_0 
       (.I0(rx_data[28]),
        .I1(TXD[28]),
        .I2(cfgRxRegData[28]),
        .O(info_o[28]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[29]_INST_0 
       (.I0(rx_data[29]),
        .I1(TXD[29]),
        .I2(cfgRxRegData[29]),
        .O(info_o[29]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[2]_INST_0 
       (.I0(rdata[2]),
        .I1(outputs[2]),
        .I2(TXD[2]),
        .I3(dat_o[2]),
        .I4(DO[2]),
        .I5(rx_data[2]),
        .O(info_o[2]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[30]_INST_0 
       (.I0(rx_data[30]),
        .I1(TXD[30]),
        .I2(cfgRxRegData[30]),
        .O(info_o[30]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[31]_INST_0 
       (.I0(rx_data[31]),
        .I1(TXD[31]),
        .I2(cfgRxRegData[31]),
        .O(info_o[31]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[3]_INST_0 
       (.I0(rdata[3]),
        .I1(outputs[3]),
        .I2(TXD[3]),
        .I3(dat_o[3]),
        .I4(DO[3]),
        .I5(rx_data[3]),
        .O(info_o[3]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[4]_INST_0 
       (.I0(rdata[4]),
        .I1(outputs[4]),
        .I2(TXD[4]),
        .I3(dat_o[4]),
        .I4(DO[4]),
        .I5(rx_data[4]),
        .O(info_o[4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[5]_INST_0 
       (.I0(rdata[5]),
        .I1(outputs[5]),
        .I2(TXD[5]),
        .I3(dat_o[5]),
        .I4(DO[5]),
        .I5(rx_data[5]),
        .O(info_o[5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[6]_INST_0 
       (.I0(rdata[6]),
        .I1(outputs[6]),
        .I2(TXD[6]),
        .I3(dat_o[6]),
        .I4(DO[6]),
        .I5(rx_data[6]),
        .O(info_o[6]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \info_o[7]_INST_0 
       (.I0(rdata[7]),
        .I1(outputs[7]),
        .I2(TXD[7]),
        .I3(dat_o[7]),
        .I4(DO[7]),
        .I5(rx_data[7]),
        .O(info_o[7]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[8]_INST_0 
       (.I0(rx_data[8]),
        .I1(DO[8]),
        .I2(rdata[8]),
        .I3(TXD[8]),
        .O(info_o[8]));
  LUT4 #(
    .INIT(16'h6996)) 
    \info_o[9]_INST_0 
       (.I0(rx_data[9]),
        .I1(DO[9]),
        .I2(rdata[9]),
        .I3(TXD[9]),
        .O(info_o[9]));
  LUT1 #(
    .INIT(2'h2)) 
    m_en_inst
       (.I0(crc_en),
        .O(m_en));
  LUT1 #(
    .INIT(2'h2)) 
    m_we_inst
       (.I0(wdata[2]),
        .O(m_we[1]));
  LUT1 #(
    .INIT(2'h2)) 
    m_we_inst__0
       (.I0(wdata[1]),
        .O(m_we[0]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst
       (.I0(inputs[3]),
        .O(mgmt_addr[9]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__0
       (.I0(inputs[2]),
        .O(mgmt_addr[8]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__1
       (.I0(inputs[1]),
        .O(mgmt_addr[7]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__2
       (.I0(inputs[0]),
        .O(mgmt_addr[6]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__3
       (.I0(mgmt_wr_data[23]),
        .O(mgmt_addr[5]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__4
       (.I0(mgmt_wr_data[22]),
        .O(mgmt_addr[4]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__5
       (.I0(mgmt_wr_data[21]),
        .O(mgmt_addr[3]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__6
       (.I0(mgmt_wr_data[20]),
        .O(mgmt_addr[2]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__7
       (.I0(mgmt_wr_data[19]),
        .O(mgmt_addr[1]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_addr_inst__8
       (.I0(mgmt_wr_data[18]),
        .O(mgmt_addr[0]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_miim_sel_inst
       (.I0(inputs[4]),
        .O(mgmt_miim_sel));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_opcode_inst
       (.I0(mgmt_wr_data[17]),
        .O(mgmt_opcode[1]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_opcode_inst__0
       (.I0(mgmt_wr_data[16]),
        .O(mgmt_opcode[0]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_req_inst
       (.I0(inputs[5]),
        .O(mgmt_req));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst
       (.I0(inputs[7]),
        .O(mgmt_wr_data[31]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__0
       (.I0(inputs[6]),
        .O(mgmt_wr_data[30]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__1
       (.I0(inputs[5]),
        .O(mgmt_wr_data[29]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__10
       (.I0(wdata[12]),
        .O(mgmt_wr_data[12]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__11
       (.I0(wdata[11]),
        .O(mgmt_wr_data[11]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__12
       (.I0(wdata[10]),
        .O(mgmt_wr_data[10]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__13
       (.I0(wdata[9]),
        .O(mgmt_wr_data[9]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__14
       (.I0(wdata[8]),
        .O(mgmt_wr_data[8]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__15
       (.I0(dat_i),
        .O(mgmt_wr_data[7]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__16
       (.I0(wdata[6]),
        .O(mgmt_wr_data[6]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__17
       (.I0(wdata[5]),
        .O(mgmt_wr_data[5]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__18
       (.I0(wdata[4]),
        .O(mgmt_wr_data[4]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__19
       (.I0(wdata[3]),
        .O(mgmt_wr_data[3]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__2
       (.I0(inputs[4]),
        .O(mgmt_wr_data[28]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__20
       (.I0(wdata[2]),
        .O(mgmt_wr_data[2]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__21
       (.I0(wdata[1]),
        .O(mgmt_wr_data[1]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__22
       (.I0(crc_en),
        .O(mgmt_wr_data[0]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__3
       (.I0(inputs[3]),
        .O(mgmt_wr_data[27]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__4
       (.I0(inputs[2]),
        .O(mgmt_wr_data[26]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__5
       (.I0(inputs[1]),
        .O(mgmt_wr_data[25]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__6
       (.I0(inputs[0]),
        .O(mgmt_wr_data[24]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__7
       (.I0(wdata[15]),
        .O(mgmt_wr_data[15]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__8
       (.I0(wdata[14]),
        .O(mgmt_wr_data[14]));
  LUT1 #(
    .INIT(2'h2)) 
    mgmt_wr_data_inst__9
       (.I0(wdata[13]),
        .O(mgmt_wr_data[13]));
  LUT1 #(
    .INIT(2'h2)) 
    miso_i_inst
       (.I0(wdata[15]),
        .O(miso_i));
  LUT1 #(
    .INIT(2'h2)) 
    run_in_inst
       (.I0(inputs[7]),
        .O(run_in));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst
       (.I0(rxStatRegPlus[6]),
        .O(dat_i_vec[6]));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst__0
       (.I0(rxStatRegPlus[5]),
        .O(dat_i_vec[5]));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst__1
       (.I0(rxStatRegPlus[4]),
        .O(dat_i_vec[4]));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst__2
       (.I0(rxStatRegPlus[3]),
        .O(dat_i_vec[3]));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst__3
       (.I0(rxStatRegPlus[2]),
        .O(dat_i_vec[2]));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst__4
       (.I0(rxStatRegPlus[1]),
        .O(dat_i_vec[1]));
  LUT1 #(
    .INIT(2'h2)) 
    rxStatRegPlus_inst__5
       (.I0(rxStatRegPlus[0]),
        .O(dat_i_vec[0]));
  LUT1 #(
    .INIT(2'h2)) 
    stb_i_inst
       (.I0(wdata[3]),
        .O(stb_i));
  LUT1 #(
    .INIT(2'h2)) 
    wdata_inst
       (.I0(dat_i),
        .O(wdata[7]));
  LUT1 #(
    .INIT(2'h2)) 
    wdata_inst__0
       (.I0(crc_en),
        .O(wdata[0]));
  LUT1 #(
    .INIT(2'h2)) 
    we_i_inst
       (.I0(wdata[6]),
        .O(we_i));
  LUT1 #(
    .INIT(2'h2)) 
    xgmii_rxc_inst
       (.I0(wdata[5]),
        .O(xgmii_rxc[3]));
  LUT1 #(
    .INIT(2'h2)) 
    xgmii_rxc_inst__0
       (.I0(wdata[4]),
        .O(xgmii_rxc[2]));
  LUT1 #(
    .INIT(2'h2)) 
    xgmii_rxc_inst__1
       (.I0(wdata[3]),
        .O(xgmii_rxc[1]));
  LUT1 #(
    .INIT(2'h2)) 
    xgmii_rxc_inst__2
       (.I0(wdata[2]),
        .O(xgmii_rxc[0]));
  LUT1 #(
    .INIT(2'h1)) 
    \xgmii_rxd[0]_i_1 
       (.I0(xgmii_rxd[0]),
        .O(\xgmii_rxd[0]_i_1_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[0] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd[0]_i_1_n_0 ),
        .Q(xgmii_rxd[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[10] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_14 ),
        .Q(xgmii_rxd[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[11] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_13 ),
        .Q(xgmii_rxd[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[12] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_12 ),
        .Q(xgmii_rxd[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[13] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_11 ),
        .Q(xgmii_rxd[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[14] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_10 ),
        .Q(xgmii_rxd[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[15] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_9 ),
        .Q(xgmii_rxd[15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[16] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_8 ),
        .Q(xgmii_rxd[16]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \xgmii_rxd_reg[16]_i_1 
       (.CI(\xgmii_rxd_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\xgmii_rxd_reg[16]_i_1_n_0 ,\xgmii_rxd_reg[16]_i_1_n_1 ,\xgmii_rxd_reg[16]_i_1_n_2 ,\xgmii_rxd_reg[16]_i_1_n_3 ,\xgmii_rxd_reg[16]_i_1_n_4 ,\xgmii_rxd_reg[16]_i_1_n_5 ,\xgmii_rxd_reg[16]_i_1_n_6 ,\xgmii_rxd_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\xgmii_rxd_reg[16]_i_1_n_8 ,\xgmii_rxd_reg[16]_i_1_n_9 ,\xgmii_rxd_reg[16]_i_1_n_10 ,\xgmii_rxd_reg[16]_i_1_n_11 ,\xgmii_rxd_reg[16]_i_1_n_12 ,\xgmii_rxd_reg[16]_i_1_n_13 ,\xgmii_rxd_reg[16]_i_1_n_14 ,\xgmii_rxd_reg[16]_i_1_n_15 }),
        .S(xgmii_rxd[16:9]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[17] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_15 ),
        .Q(xgmii_rxd[17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[18] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_14 ),
        .Q(xgmii_rxd[18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[19] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_13 ),
        .Q(xgmii_rxd[19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[1] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_15 ),
        .Q(xgmii_rxd[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[20] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_12 ),
        .Q(xgmii_rxd[20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[21] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_11 ),
        .Q(xgmii_rxd[21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[22] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_10 ),
        .Q(xgmii_rxd[22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[23] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_9 ),
        .Q(xgmii_rxd[23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[24] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[24]_i_1_n_8 ),
        .Q(xgmii_rxd[24]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \xgmii_rxd_reg[24]_i_1 
       (.CI(\xgmii_rxd_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\xgmii_rxd_reg[24]_i_1_n_0 ,\xgmii_rxd_reg[24]_i_1_n_1 ,\xgmii_rxd_reg[24]_i_1_n_2 ,\xgmii_rxd_reg[24]_i_1_n_3 ,\xgmii_rxd_reg[24]_i_1_n_4 ,\xgmii_rxd_reg[24]_i_1_n_5 ,\xgmii_rxd_reg[24]_i_1_n_6 ,\xgmii_rxd_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\xgmii_rxd_reg[24]_i_1_n_8 ,\xgmii_rxd_reg[24]_i_1_n_9 ,\xgmii_rxd_reg[24]_i_1_n_10 ,\xgmii_rxd_reg[24]_i_1_n_11 ,\xgmii_rxd_reg[24]_i_1_n_12 ,\xgmii_rxd_reg[24]_i_1_n_13 ,\xgmii_rxd_reg[24]_i_1_n_14 ,\xgmii_rxd_reg[24]_i_1_n_15 }),
        .S(xgmii_rxd[24:17]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[25] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_15 ),
        .Q(xgmii_rxd[25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[26] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_14 ),
        .Q(xgmii_rxd[26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[27] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_13 ),
        .Q(xgmii_rxd[27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[28] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_12 ),
        .Q(xgmii_rxd[28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[29] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_11 ),
        .Q(xgmii_rxd[29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[2] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_14 ),
        .Q(xgmii_rxd[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[30] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_10 ),
        .Q(xgmii_rxd[30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[31] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[31]_i_1_n_9 ),
        .Q(xgmii_rxd[31]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \xgmii_rxd_reg[31]_i_1 
       (.CI(\xgmii_rxd_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_xgmii_rxd_reg[31]_i_1_CO_UNCONNECTED [7:6],\xgmii_rxd_reg[31]_i_1_n_2 ,\xgmii_rxd_reg[31]_i_1_n_3 ,\xgmii_rxd_reg[31]_i_1_n_4 ,\xgmii_rxd_reg[31]_i_1_n_5 ,\xgmii_rxd_reg[31]_i_1_n_6 ,\xgmii_rxd_reg[31]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_xgmii_rxd_reg[31]_i_1_O_UNCONNECTED [7],\xgmii_rxd_reg[31]_i_1_n_9 ,\xgmii_rxd_reg[31]_i_1_n_10 ,\xgmii_rxd_reg[31]_i_1_n_11 ,\xgmii_rxd_reg[31]_i_1_n_12 ,\xgmii_rxd_reg[31]_i_1_n_13 ,\xgmii_rxd_reg[31]_i_1_n_14 ,\xgmii_rxd_reg[31]_i_1_n_15 }),
        .S({1'b0,xgmii_rxd[31:25]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[3] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_13 ),
        .Q(xgmii_rxd[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[4] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_12 ),
        .Q(xgmii_rxd[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[5] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_11 ),
        .Q(xgmii_rxd[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[6] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_10 ),
        .Q(xgmii_rxd[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[7] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_9 ),
        .Q(xgmii_rxd[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[8] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[8]_i_1_n_8 ),
        .Q(xgmii_rxd[8]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \xgmii_rxd_reg[8]_i_1 
       (.CI(xgmii_rxd[0]),
        .CI_TOP(1'b0),
        .CO({\xgmii_rxd_reg[8]_i_1_n_0 ,\xgmii_rxd_reg[8]_i_1_n_1 ,\xgmii_rxd_reg[8]_i_1_n_2 ,\xgmii_rxd_reg[8]_i_1_n_3 ,\xgmii_rxd_reg[8]_i_1_n_4 ,\xgmii_rxd_reg[8]_i_1_n_5 ,\xgmii_rxd_reg[8]_i_1_n_6 ,\xgmii_rxd_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\xgmii_rxd_reg[8]_i_1_n_8 ,\xgmii_rxd_reg[8]_i_1_n_9 ,\xgmii_rxd_reg[8]_i_1_n_10 ,\xgmii_rxd_reg[8]_i_1_n_11 ,\xgmii_rxd_reg[8]_i_1_n_12 ,\xgmii_rxd_reg[8]_i_1_n_13 ,\xgmii_rxd_reg[8]_i_1_n_14 ,\xgmii_rxd_reg[8]_i_1_n_15 }),
        .S(xgmii_rxd[8:1]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \xgmii_rxd_reg[9] 
       (.C(rxclk_out),
        .CE(1'b1),
        .D(\xgmii_rxd_reg[16]_i_1_n_15 ),
        .Q(xgmii_rxd[9]),
        .R(1'b0));
endmodule

(* ORIG_REF_NAME = "CRC32_D64" *) 
module switch_elements_CRC32_D64
   (Q,
    frame_start_del,
    transmit_pause_frame_valid,
    SS,
    clk_i,
    \CRC_OUT_reg[24]_0 );
  output [31:0]Q;
  input frame_start_del;
  input transmit_pause_frame_valid;
  input [0:0]SS;
  input clk_i;
  input [63:0]\CRC_OUT_reg[24]_0 ;

  wire \CRC_OUT[0]_i_2__0_n_0 ;
  wire \CRC_OUT[0]_i_3__0_n_0 ;
  wire \CRC_OUT[0]_i_4__0_n_0 ;
  wire \CRC_OUT[10]_i_2__1_n_0 ;
  wire \CRC_OUT[10]_i_3__1_n_0 ;
  wire \CRC_OUT[10]_i_4__0_n_0 ;
  wire \CRC_OUT[10]_i_5__0_n_0 ;
  wire \CRC_OUT[11]_i_2__1_n_0 ;
  wire \CRC_OUT[11]_i_3__0_n_0 ;
  wire \CRC_OUT[11]_i_4__0_n_0 ;
  wire \CRC_OUT[11]_i_5__0_n_0 ;
  wire \CRC_OUT[11]_i_6__0_n_0 ;
  wire \CRC_OUT[12]_i_2__1_n_0 ;
  wire \CRC_OUT[12]_i_3__0_n_0 ;
  wire \CRC_OUT[12]_i_4__0_n_0 ;
  wire \CRC_OUT[12]_i_5__0_n_0 ;
  wire \CRC_OUT[12]_i_6__0_n_0 ;
  wire \CRC_OUT[13]_i_2__1_n_0 ;
  wire \CRC_OUT[13]_i_3__1_n_0 ;
  wire \CRC_OUT[13]_i_4__0_n_0 ;
  wire \CRC_OUT[13]_i_5__0_n_0 ;
  wire \CRC_OUT[13]_i_6__0_n_0 ;
  wire \CRC_OUT[13]_i_7__0_n_0 ;
  wire \CRC_OUT[14]_i_2__0_n_0 ;
  wire \CRC_OUT[14]_i_3__1_n_0 ;
  wire \CRC_OUT[14]_i_4__0_n_0 ;
  wire \CRC_OUT[14]_i_5__0_n_0 ;
  wire \CRC_OUT[15]_i_2__1_n_0 ;
  wire \CRC_OUT[15]_i_3__1_n_0 ;
  wire \CRC_OUT[15]_i_4__0_n_0 ;
  wire \CRC_OUT[16]_i_2__1_n_0 ;
  wire \CRC_OUT[16]_i_3__1_n_0 ;
  wire \CRC_OUT[16]_i_4__1_n_0 ;
  wire \CRC_OUT[16]_i_5__0_n_0 ;
  wire \CRC_OUT[17]_i_2__1_n_0 ;
  wire \CRC_OUT[17]_i_3__0_n_0 ;
  wire \CRC_OUT[17]_i_4__0_n_0 ;
  wire \CRC_OUT[17]_i_5__0_n_0 ;
  wire \CRC_OUT[17]_i_6__0_n_0 ;
  wire \CRC_OUT[17]_i_7__0_n_0 ;
  wire \CRC_OUT[17]_i_8__0_n_0 ;
  wire \CRC_OUT[18]_i_2__0_n_0 ;
  wire \CRC_OUT[18]_i_3__1_n_0 ;
  wire \CRC_OUT[18]_i_4__0_n_0 ;
  wire \CRC_OUT[18]_i_5__0_n_0 ;
  wire \CRC_OUT[18]_i_6__0_n_0 ;
  wire \CRC_OUT[18]_i_7__0_n_0 ;
  wire \CRC_OUT[19]_i_2__1_n_0 ;
  wire \CRC_OUT[19]_i_3__0_n_0 ;
  wire \CRC_OUT[19]_i_4__0_n_0 ;
  wire \CRC_OUT[19]_i_5__0_n_0 ;
  wire \CRC_OUT[19]_i_6__0_n_0 ;
  wire \CRC_OUT[1]_i_2__0_n_0 ;
  wire \CRC_OUT[1]_i_3__0_n_0 ;
  wire \CRC_OUT[1]_i_4__0_n_0 ;
  wire \CRC_OUT[20]_i_2__0_n_0 ;
  wire \CRC_OUT[20]_i_3__0_n_0 ;
  wire \CRC_OUT[20]_i_4__0_n_0 ;
  wire \CRC_OUT[20]_i_5__0_n_0 ;
  wire \CRC_OUT[21]_i_2__0_n_0 ;
  wire \CRC_OUT[21]_i_3__0_n_0 ;
  wire \CRC_OUT[21]_i_4__0_n_0 ;
  wire \CRC_OUT[22]_i_2__0_n_0 ;
  wire \CRC_OUT[22]_i_3__0_n_0 ;
  wire \CRC_OUT[22]_i_4__0_n_0 ;
  wire \CRC_OUT[22]_i_5__0_n_0 ;
  wire \CRC_OUT[22]_i_6__0_n_0 ;
  wire \CRC_OUT[22]_i_7__0_n_0 ;
  wire \CRC_OUT[23]_i_2__1_n_0 ;
  wire \CRC_OUT[23]_i_3__0_n_0 ;
  wire \CRC_OUT[23]_i_4__0_n_0 ;
  wire \CRC_OUT[23]_i_5__0_n_0 ;
  wire \CRC_OUT[23]_i_6__0_n_0 ;
  wire \CRC_OUT[23]_i_7__0_n_0 ;
  wire \CRC_OUT[23]_i_8__0_n_0 ;
  wire \CRC_OUT[24]_i_10__0_n_0 ;
  wire \CRC_OUT[24]_i_11__0_n_0 ;
  wire \CRC_OUT[24]_i_12__0_n_0 ;
  wire \CRC_OUT[24]_i_2__1_n_0 ;
  wire \CRC_OUT[24]_i_3__1_n_0 ;
  wire \CRC_OUT[24]_i_4__1_n_0 ;
  wire \CRC_OUT[24]_i_5__0_n_0 ;
  wire \CRC_OUT[24]_i_6__0_n_0 ;
  wire \CRC_OUT[24]_i_7__0_n_0 ;
  wire \CRC_OUT[24]_i_8__0_n_0 ;
  wire \CRC_OUT[24]_i_9__0_n_0 ;
  wire \CRC_OUT[25]_i_10__0_n_0 ;
  wire \CRC_OUT[25]_i_2__1_n_0 ;
  wire \CRC_OUT[25]_i_3__0_n_0 ;
  wire \CRC_OUT[25]_i_4__0_n_0 ;
  wire \CRC_OUT[25]_i_5__0_n_0 ;
  wire \CRC_OUT[25]_i_6__0_n_0 ;
  wire \CRC_OUT[25]_i_7__0_n_0 ;
  wire \CRC_OUT[25]_i_8__0_n_0 ;
  wire \CRC_OUT[25]_i_9__0_n_0 ;
  wire \CRC_OUT[26]_i_2__1_n_0 ;
  wire \CRC_OUT[26]_i_3__0_n_0 ;
  wire \CRC_OUT[26]_i_4__0_n_0 ;
  wire \CRC_OUT[26]_i_5__0_n_0 ;
  wire \CRC_OUT[26]_i_6__0_n_0 ;
  wire \CRC_OUT[26]_i_7__0_n_0 ;
  wire \CRC_OUT[26]_i_8__0_n_0 ;
  wire \CRC_OUT[27]_i_2__1_n_0 ;
  wire \CRC_OUT[27]_i_3__0_n_0 ;
  wire \CRC_OUT[27]_i_4__0_n_0 ;
  wire \CRC_OUT[27]_i_5__0_n_0 ;
  wire \CRC_OUT[27]_i_6__0_n_0 ;
  wire \CRC_OUT[27]_i_7__0_n_0 ;
  wire \CRC_OUT[27]_i_8__0_n_0 ;
  wire \CRC_OUT[28]_i_10__0_n_0 ;
  wire \CRC_OUT[28]_i_11__0_n_0 ;
  wire \CRC_OUT[28]_i_12__0_n_0 ;
  wire \CRC_OUT[28]_i_2__1_n_0 ;
  wire \CRC_OUT[28]_i_3__0_n_0 ;
  wire \CRC_OUT[28]_i_4__0_n_0 ;
  wire \CRC_OUT[28]_i_5__0_n_0 ;
  wire \CRC_OUT[28]_i_6__0_n_0 ;
  wire \CRC_OUT[28]_i_7__0_n_0 ;
  wire \CRC_OUT[28]_i_8__0_n_0 ;
  wire \CRC_OUT[28]_i_9__0_n_0 ;
  wire \CRC_OUT[29]_i_2__1_n_0 ;
  wire \CRC_OUT[29]_i_3__0_n_0 ;
  wire \CRC_OUT[29]_i_4__0_n_0 ;
  wire \CRC_OUT[29]_i_5__0_n_0 ;
  wire \CRC_OUT[29]_i_6__0_n_0 ;
  wire \CRC_OUT[29]_i_7__0_n_0 ;
  wire \CRC_OUT[29]_i_8__0_n_0 ;
  wire \CRC_OUT[2]_i_2__1_n_0 ;
  wire \CRC_OUT[2]_i_3__0_n_0 ;
  wire \CRC_OUT[2]_i_4__0_n_0 ;
  wire \CRC_OUT[2]_i_5__0_n_0 ;
  wire \CRC_OUT[30]_i_10__0_n_0 ;
  wire \CRC_OUT[30]_i_11__0_n_0 ;
  wire \CRC_OUT[30]_i_2__1_n_0 ;
  wire \CRC_OUT[30]_i_3__0_n_0 ;
  wire \CRC_OUT[30]_i_4__0_n_0 ;
  wire \CRC_OUT[30]_i_5__0_n_0 ;
  wire \CRC_OUT[30]_i_6__0_n_0 ;
  wire \CRC_OUT[30]_i_7__0_n_0 ;
  wire \CRC_OUT[30]_i_8__0_n_0 ;
  wire \CRC_OUT[30]_i_9__0_n_0 ;
  wire \CRC_OUT[31]_i_10__0_n_0 ;
  wire \CRC_OUT[31]_i_11__0_n_0 ;
  wire \CRC_OUT[31]_i_12_n_0 ;
  wire \CRC_OUT[31]_i_2__0_n_0 ;
  wire \CRC_OUT[31]_i_4__0_n_0 ;
  wire \CRC_OUT[31]_i_5__0_n_0 ;
  wire \CRC_OUT[31]_i_6__0_n_0 ;
  wire \CRC_OUT[31]_i_7__0_n_0 ;
  wire \CRC_OUT[31]_i_8__0_n_0 ;
  wire \CRC_OUT[31]_i_9__0_n_0 ;
  wire \CRC_OUT[3]_i_2__0_n_0 ;
  wire \CRC_OUT[3]_i_3__0_n_0 ;
  wire \CRC_OUT[4]_i_2__1_n_0 ;
  wire \CRC_OUT[4]_i_3__0_n_0 ;
  wire \CRC_OUT[4]_i_4__0_n_0 ;
  wire \CRC_OUT[5]_i_2__1_n_0 ;
  wire \CRC_OUT[5]_i_3__0_n_0 ;
  wire \CRC_OUT[5]_i_4__0_n_0 ;
  wire \CRC_OUT[5]_i_5__0_n_0 ;
  wire \CRC_OUT[5]_i_6__0_n_0 ;
  wire \CRC_OUT[6]_i_2__1_n_0 ;
  wire \CRC_OUT[6]_i_3__0_n_0 ;
  wire \CRC_OUT[7]_i_2__1_n_0 ;
  wire \CRC_OUT[7]_i_3__0_n_0 ;
  wire \CRC_OUT[7]_i_4__0_n_0 ;
  wire \CRC_OUT[7]_i_5__0_n_0 ;
  wire \CRC_OUT[8]_i_2__0_n_0 ;
  wire \CRC_OUT[8]_i_3__0_n_0 ;
  wire \CRC_OUT[8]_i_4__0_n_0 ;
  wire \CRC_OUT[8]_i_5__0_n_0 ;
  wire \CRC_OUT[8]_i_6__0_n_0 ;
  wire \CRC_OUT[9]_i_2__1_n_0 ;
  wire \CRC_OUT[9]_i_3__0_n_0 ;
  wire \CRC_OUT[9]_i_4__0_n_0 ;
  wire \CRC_OUT[9]_i_5__0_n_0 ;
  wire \CRC_OUT[9]_i_6__0_n_0 ;
  wire [63:0]\CRC_OUT_reg[24]_0 ;
  wire [31:0]Q;
  wire [0:0]SS;
  wire clk_i;
  wire frame_start_del;
  wire nextCRC32_D64_return0;
  wire nextCRC32_D64_return0100_out;
  wire nextCRC32_D64_return0102_out;
  wire nextCRC32_D64_return0104_out;
  wire nextCRC32_D64_return0106_out;
  wire nextCRC32_D64_return0108_out;
  wire nextCRC32_D64_return0109_out;
  wire nextCRC32_D64_return0110_out;
  wire nextCRC32_D64_return0112_out;
  wire nextCRC32_D64_return0114_out;
  wire nextCRC32_D64_return0116_out;
  wire nextCRC32_D64_return0118_out;
  wire nextCRC32_D64_return0120_out;
  wire nextCRC32_D64_return0122_out;
  wire nextCRC32_D64_return0124_out;
  wire nextCRC32_D64_return0126_out;
  wire nextCRC32_D64_return0128_out;
  wire nextCRC32_D64_return0130_out;
  wire nextCRC32_D64_return0132_out;
  wire nextCRC32_D64_return0134_out;
  wire nextCRC32_D64_return0136_out;
  wire nextCRC32_D64_return0138_out;
  wire nextCRC32_D64_return056_out;
  wire nextCRC32_D64_return068_out;
  wire nextCRC32_D64_return075_out;
  wire nextCRC32_D64_return080_out;
  wire nextCRC32_D64_return086_out;
  wire nextCRC32_D64_return091_out;
  wire nextCRC32_D64_return093_out;
  wire nextCRC32_D64_return094_out;
  wire nextCRC32_D64_return096_out;
  wire nextCRC32_D64_return098_out;
  wire transmit_pause_frame_valid;

  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[0]_i_1__1 
       (.I0(\CRC_OUT[0]_i_2__0_n_0 ),
        .I1(\CRC_OUT[20]_i_2__0_n_0 ),
        .I2(\CRC_OUT[12]_i_2__1_n_0 ),
        .I3(\CRC_OUT[0]_i_3__0_n_0 ),
        .I4(\CRC_OUT[27]_i_3__0_n_0 ),
        .I5(\CRC_OUT[0]_i_4__0_n_0 ),
        .O(nextCRC32_D64_return0));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[0]_i_2__0 
       (.I0(\CRC_OUT[10]_i_3__1_n_0 ),
        .I1(\CRC_OUT[22]_i_6__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [6]),
        .I3(\CRC_OUT_reg[24]_0 [0]),
        .I4(\CRC_OUT[31]_i_12_n_0 ),
        .I5(\CRC_OUT[13]_i_7__0_n_0 ),
        .O(\CRC_OUT[0]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[0]_i_3__0 
       (.I0(\CRC_OUT_reg[24]_0 [30]),
        .I1(\CRC_OUT_reg[24]_0 [28]),
        .O(\CRC_OUT[0]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair358" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[0]_i_4__0 
       (.I0(\CRC_OUT[7]_i_4__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [29]),
        .I2(Q[15]),
        .I3(\CRC_OUT_reg[24]_0 [47]),
        .O(\CRC_OUT[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[10]_i_1__1 
       (.I0(\CRC_OUT[10]_i_2__1_n_0 ),
        .I1(\CRC_OUT[10]_i_3__1_n_0 ),
        .I2(\CRC_OUT[10]_i_4__0_n_0 ),
        .I3(\CRC_OUT[10]_i_5__0_n_0 ),
        .I4(\CRC_OUT[11]_i_6__0_n_0 ),
        .I5(\CRC_OUT[27]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return098_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[10]_i_2__1 
       (.I0(Q[24]),
        .I1(\CRC_OUT_reg[24]_0 [56]),
        .I2(\CRC_OUT[17]_i_8__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [2]),
        .I4(Q[20]),
        .I5(\CRC_OUT_reg[24]_0 [52]),
        .O(\CRC_OUT[10]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair363" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[10]_i_3__1 
       (.I0(\CRC_OUT_reg[24]_0 [32]),
        .I1(Q[0]),
        .I2(\CRC_OUT_reg[24]_0 [58]),
        .I3(Q[26]),
        .O(\CRC_OUT[10]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair355" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[10]_i_4__0 
       (.I0(Q[30]),
        .I1(\CRC_OUT_reg[24]_0 [62]),
        .O(\CRC_OUT[10]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair340" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[10]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [13]),
        .I1(\CRC_OUT_reg[24]_0 [5]),
        .I2(\CRC_OUT[30]_i_7__0_n_0 ),
        .I3(\CRC_OUT[19]_i_4__0_n_0 ),
        .I4(\CRC_OUT[26]_i_2__1_n_0 ),
        .O(\CRC_OUT[10]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_1__1 
       (.I0(\CRC_OUT[11]_i_2__1_n_0 ),
        .I1(\CRC_OUT[11]_i_3__0_n_0 ),
        .I2(\CRC_OUT[11]_i_4__0_n_0 ),
        .I3(\CRC_OUT[11]_i_5__0_n_0 ),
        .I4(\CRC_OUT[11]_i_6__0_n_0 ),
        .I5(\CRC_OUT[29]_i_7__0_n_0 ),
        .O(nextCRC32_D64_return0100_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_2__1 
       (.I0(Q[8]),
        .I1(\CRC_OUT_reg[24]_0 [40]),
        .I2(\CRC_OUT_reg[24]_0 [43]),
        .I3(Q[11]),
        .I4(\CRC_OUT_reg[24]_0 [16]),
        .I5(\CRC_OUT[17]_i_8__0_n_0 ),
        .O(\CRC_OUT[11]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair371" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[11]_i_3__0 
       (.I0(\CRC_OUT_reg[24]_0 [20]),
        .I1(\CRC_OUT_reg[24]_0 [4]),
        .O(\CRC_OUT[11]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair365" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[11]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [3]),
        .I1(\CRC_OUT_reg[24]_0 [28]),
        .O(\CRC_OUT[11]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_5__0 
       (.I0(\CRC_OUT[28]_i_4__0_n_0 ),
        .I1(Q[16]),
        .I2(\CRC_OUT_reg[24]_0 [48]),
        .I3(\CRC_OUT[28]_i_9__0_n_0 ),
        .I4(\CRC_OUT[31]_i_4__0_n_0 ),
        .I5(\CRC_OUT[24]_i_2__1_n_0 ),
        .O(\CRC_OUT[11]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair333" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[11]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [0]),
        .I1(\CRC_OUT[22]_i_5__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [26]),
        .I3(Q[23]),
        .I4(\CRC_OUT_reg[24]_0 [55]),
        .O(\CRC_OUT[11]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[12]_i_1__1 
       (.I0(\CRC_OUT[20]_i_4__0_n_0 ),
        .I1(\CRC_OUT[12]_i_2__1_n_0 ),
        .I2(\CRC_OUT[12]_i_3__0_n_0 ),
        .I3(\CRC_OUT[12]_i_4__0_n_0 ),
        .I4(\CRC_OUT[23]_i_5__0_n_0 ),
        .I5(\CRC_OUT[12]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0102_out));
  (* SOFT_HLUTNM = "soft_lutpair354" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[12]_i_2__1 
       (.I0(\CRC_OUT_reg[24]_0 [31]),
        .I1(\CRC_OUT_reg[24]_0 [9]),
        .I2(\CRC_OUT_reg[24]_0 [63]),
        .I3(Q[31]),
        .O(\CRC_OUT[12]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[12]_i_3__0 
       (.I0(\CRC_OUT[31]_i_4__0_n_0 ),
        .I1(\CRC_OUT[26]_i_3__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [18]),
        .I3(\CRC_OUT_reg[24]_0 [2]),
        .I4(\CRC_OUT_reg[24]_0 [5]),
        .I5(\CRC_OUT_reg[24]_0 [21]),
        .O(\CRC_OUT[12]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[12]_i_4__0 
       (.I0(\CRC_OUT[12]_i_6__0_n_0 ),
        .I1(\CRC_OUT[30]_i_11__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [30]),
        .I3(\CRC_OUT_reg[24]_0 [24]),
        .I4(\CRC_OUT[28]_i_12__0_n_0 ),
        .I5(\CRC_OUT[28]_i_9__0_n_0 ),
        .O(\CRC_OUT[12]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair359" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[12]_i_5__0 
       (.I0(Q[29]),
        .I1(\CRC_OUT_reg[24]_0 [61]),
        .I2(Q[21]),
        .I3(\CRC_OUT_reg[24]_0 [53]),
        .O(\CRC_OUT[12]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair346" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[12]_i_6__0 
       (.I0(Q[10]),
        .I1(\CRC_OUT_reg[24]_0 [42]),
        .O(\CRC_OUT[12]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_1__1 
       (.I0(\CRC_OUT[13]_i_2__1_n_0 ),
        .I1(\CRC_OUT[13]_i_3__1_n_0 ),
        .I2(\CRC_OUT[13]_i_4__0_n_0 ),
        .I3(\CRC_OUT[13]_i_5__0_n_0 ),
        .I4(\CRC_OUT[30]_i_5__0_n_0 ),
        .I5(\CRC_OUT[13]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return0104_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_2__1 
       (.I0(\CRC_OUT[10]_i_4__0_n_0 ),
        .I1(\CRC_OUT[24]_i_12__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [5]),
        .I3(\CRC_OUT_reg[24]_0 [25]),
        .I4(\CRC_OUT[13]_i_7__0_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 [10]),
        .O(\CRC_OUT[13]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_3__1 
       (.I0(\CRC_OUT_reg[24]_0 [6]),
        .I1(\CRC_OUT_reg[24]_0 [13]),
        .I2(\CRC_OUT_reg[24]_0 [18]),
        .I3(\CRC_OUT_reg[24]_0 [2]),
        .I4(\CRC_OUT[19]_i_4__0_n_0 ),
        .I5(\CRC_OUT[11]_i_4__0_n_0 ),
        .O(\CRC_OUT[13]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair366" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[13]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [55]),
        .I1(Q[23]),
        .I2(\CRC_OUT_reg[24]_0 [1]),
        .O(\CRC_OUT[13]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair347" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[13]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [22]),
        .I1(Q[10]),
        .I2(\CRC_OUT_reg[24]_0 [42]),
        .I3(\CRC_OUT[30]_i_11__0_n_0 ),
        .O(\CRC_OUT[13]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair335" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[13]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [31]),
        .I1(\CRC_OUT_reg[24]_0 [19]),
        .I2(\CRC_OUT_reg[24]_0 [48]),
        .I3(Q[16]),
        .I4(\CRC_OUT[31]_i_11__0_n_0 ),
        .O(\CRC_OUT[13]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair350" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[13]_i_7__0 
       (.I0(Q[22]),
        .I1(\CRC_OUT_reg[24]_0 [54]),
        .O(\CRC_OUT[13]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[14]_i_1__1 
       (.I0(\CRC_OUT[14]_i_2__0_n_0 ),
        .I1(\CRC_OUT[19]_i_5__0_n_0 ),
        .I2(\CRC_OUT[30]_i_5__0_n_0 ),
        .I3(\CRC_OUT[27]_i_3__0_n_0 ),
        .I4(\CRC_OUT[14]_i_3__1_n_0 ),
        .I5(\CRC_OUT[14]_i_4__0_n_0 ),
        .O(nextCRC32_D64_return0106_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[14]_i_2__0 
       (.I0(\CRC_OUT[14]_i_5__0_n_0 ),
        .I1(\CRC_OUT[11]_i_3__0_n_0 ),
        .I2(\CRC_OUT[28]_i_12__0_n_0 ),
        .I3(\CRC_OUT[25]_i_8__0_n_0 ),
        .I4(\CRC_OUT[30]_i_11__0_n_0 ),
        .I5(\CRC_OUT[30]_i_10__0_n_0 ),
        .O(\CRC_OUT[14]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair370" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[14]_i_3__1 
       (.I0(\CRC_OUT_reg[24]_0 [6]),
        .I1(\CRC_OUT_reg[24]_0 [2]),
        .O(\CRC_OUT[14]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[14]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [11]),
        .I1(\CRC_OUT[24]_i_12__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [23]),
        .I3(\CRC_OUT_reg[24]_0 [17]),
        .I4(Q[24]),
        .I5(\CRC_OUT_reg[24]_0 [56]),
        .O(\CRC_OUT[14]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair360" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[14]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [19]),
        .I1(\CRC_OUT_reg[24]_0 [29]),
        .O(\CRC_OUT[14]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[15]_i_1__1 
       (.I0(\CRC_OUT[15]_i_2__1_n_0 ),
        .I1(\CRC_OUT[20]_i_2__0_n_0 ),
        .I2(\CRC_OUT[15]_i_3__1_n_0 ),
        .I3(\CRC_OUT[19]_i_5__0_n_0 ),
        .I4(\CRC_OUT[28]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0108_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[15]_i_2__1 
       (.I0(\CRC_OUT[24]_i_9__0_n_0 ),
        .I1(\CRC_OUT[15]_i_4__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [18]),
        .I3(\CRC_OUT_reg[24]_0 [9]),
        .I4(\CRC_OUT[17]_i_7__0_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 [30]),
        .O(\CRC_OUT[15]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[15]_i_3__1 
       (.I0(\CRC_OUT[22]_i_6__0_n_0 ),
        .I1(\CRC_OUT[27]_i_2__1_n_0 ),
        .I2(Q[13]),
        .I3(\CRC_OUT_reg[24]_0 [45]),
        .I4(\CRC_OUT[27]_i_7__0_n_0 ),
        .O(\CRC_OUT[15]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair357" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[15]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [57]),
        .I1(Q[25]),
        .O(\CRC_OUT[15]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[16]_i_1__1 
       (.I0(\CRC_OUT[16]_i_2__1_n_0 ),
        .I1(\CRC_OUT[16]_i_3__1_n_0 ),
        .I2(\CRC_OUT[17]_i_5__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [17]),
        .I4(Q[24]),
        .I5(\CRC_OUT_reg[24]_0 [56]),
        .O(nextCRC32_D64_return0109_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[16]_i_2__1 
       (.I0(\CRC_OUT[16]_i_4__1_n_0 ),
        .I1(\CRC_OUT[16]_i_5__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [4]),
        .I3(\CRC_OUT_reg[24]_0 [22]),
        .I4(\CRC_OUT_reg[24]_0 [13]),
        .I5(\CRC_OUT_reg[24]_0 [26]),
        .O(\CRC_OUT[16]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[16]_i_3__1 
       (.I0(\CRC_OUT[22]_i_4__0_n_0 ),
        .I1(\CRC_OUT[24]_i_7__0_n_0 ),
        .I2(\CRC_OUT[28]_i_4__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [30]),
        .I4(\CRC_OUT_reg[24]_0 [8]),
        .O(\CRC_OUT[16]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair364" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[16]_i_4__1 
       (.I0(\CRC_OUT_reg[24]_0 [5]),
        .I1(\CRC_OUT_reg[24]_0 [21]),
        .O(\CRC_OUT[16]_i_4__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair334" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[16]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [46]),
        .I1(Q[14]),
        .I2(\CRC_OUT_reg[24]_0 [0]),
        .O(\CRC_OUT[16]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_1__1 
       (.I0(\CRC_OUT[17]_i_2__1_n_0 ),
        .I1(\CRC_OUT[17]_i_3__0_n_0 ),
        .I2(\CRC_OUT[17]_i_4__0_n_0 ),
        .I3(\CRC_OUT[17]_i_5__0_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [20]),
        .I5(\CRC_OUT_reg[24]_0 [22]),
        .O(nextCRC32_D64_return0110_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_2__1 
       (.I0(\CRC_OUT_reg[24]_0 [18]),
        .I1(\CRC_OUT_reg[24]_0 [30]),
        .I2(\CRC_OUT_reg[24]_0 [23]),
        .I3(\CRC_OUT_reg[24]_0 [5]),
        .I4(\CRC_OUT_reg[24]_0 [27]),
        .I5(\CRC_OUT_reg[24]_0 [1]),
        .O(\CRC_OUT[17]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_3__0 
       (.I0(\CRC_OUT[17]_i_6__0_n_0 ),
        .I1(\CRC_OUT[22]_i_5__0_n_0 ),
        .I2(\CRC_OUT[28]_i_12__0_n_0 ),
        .I3(\CRC_OUT[17]_i_7__0_n_0 ),
        .I4(\CRC_OUT[26]_i_7__0_n_0 ),
        .I5(\CRC_OUT[17]_i_8__0_n_0 ),
        .O(\CRC_OUT[17]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair336" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[17]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [25]),
        .I1(Q[13]),
        .I2(\CRC_OUT_reg[24]_0 [45]),
        .I3(\CRC_OUT_reg[24]_0 [58]),
        .I4(Q[26]),
        .O(\CRC_OUT[17]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_5__0 
       (.I0(Q[15]),
        .I1(\CRC_OUT_reg[24]_0 [47]),
        .I2(\CRC_OUT_reg[24]_0 [57]),
        .I3(Q[25]),
        .I4(Q[16]),
        .I5(\CRC_OUT_reg[24]_0 [48]),
        .O(\CRC_OUT[17]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair370" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [6]),
        .I1(\CRC_OUT_reg[24]_0 [13]),
        .O(\CRC_OUT[17]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_7__0 
       (.I0(Q[20]),
        .I1(\CRC_OUT_reg[24]_0 [52]),
        .O(\CRC_OUT[17]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair343" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [33]),
        .I1(Q[1]),
        .O(\CRC_OUT[17]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[18]_i_1__1 
       (.I0(\CRC_OUT[26]_i_5__0_n_0 ),
        .I1(\CRC_OUT[18]_i_2__0_n_0 ),
        .I2(\CRC_OUT[18]_i_3__1_n_0 ),
        .I3(\CRC_OUT[18]_i_4__0_n_0 ),
        .I4(\CRC_OUT[18]_i_5__0_n_0 ),
        .I5(\CRC_OUT[20]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0112_out));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_2__0 
       (.I0(\CRC_OUT_reg[24]_0 [26]),
        .I1(\CRC_OUT_reg[24]_0 [24]),
        .O(\CRC_OUT[18]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[18]_i_3__1 
       (.I0(\CRC_OUT[14]_i_3__1_n_0 ),
        .I1(\CRC_OUT[10]_i_3__1_n_0 ),
        .I2(\CRC_OUT[27]_i_7__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [14]),
        .I4(\CRC_OUT[29]_i_4__0_n_0 ),
        .I5(\CRC_OUT[24]_i_10__0_n_0 ),
        .O(\CRC_OUT[18]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[18]_i_4__0 
       (.I0(\CRC_OUT[18]_i_6__0_n_0 ),
        .I1(\CRC_OUT[23]_i_8__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [15]),
        .I3(\CRC_OUT_reg[24]_0 [28]),
        .I4(\CRC_OUT[28]_i_12__0_n_0 ),
        .I5(\CRC_OUT[18]_i_7__0_n_0 ),
        .O(\CRC_OUT[18]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair367" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[18]_i_5__0 
       (.I0(Q[16]),
        .I1(\CRC_OUT_reg[24]_0 [48]),
        .I2(\CRC_OUT_reg[24]_0 [50]),
        .I3(Q[18]),
        .O(\CRC_OUT[18]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_6__0 
       (.I0(Q[14]),
        .I1(\CRC_OUT_reg[24]_0 [46]),
        .O(\CRC_OUT[18]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair351" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_7__0 
       (.I0(Q[27]),
        .I1(\CRC_OUT_reg[24]_0 [59]),
        .O(\CRC_OUT[18]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[19]_i_1__1 
       (.I0(\CRC_OUT[19]_i_2__1_n_0 ),
        .I1(\CRC_OUT[19]_i_3__0_n_0 ),
        .I2(\CRC_OUT[19]_i_4__0_n_0 ),
        .I3(\CRC_OUT[19]_i_5__0_n_0 ),
        .I4(\CRC_OUT[25]_i_4__0_n_0 ),
        .I5(\CRC_OUT[19]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return0114_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[19]_i_2__1 
       (.I0(\CRC_OUT[24]_i_8__0_n_0 ),
        .I1(\CRC_OUT[28]_i_12__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [7]),
        .I3(\CRC_OUT_reg[24]_0 [25]),
        .I4(\CRC_OUT_reg[24]_0 [27]),
        .I5(\CRC_OUT_reg[24]_0 [24]),
        .O(\CRC_OUT[19]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[19]_i_3__0 
       (.I0(Q[0]),
        .I1(\CRC_OUT_reg[24]_0 [32]),
        .I2(\CRC_OUT_reg[24]_0 [35]),
        .I3(Q[3]),
        .I4(\CRC_OUT_reg[24]_0 [22]),
        .I5(\CRC_OUT_reg[24]_0 [20]),
        .O(\CRC_OUT[19]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair349" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[19]_i_4__0 
       (.I0(Q[18]),
        .I1(\CRC_OUT_reg[24]_0 [50]),
        .I2(\CRC_OUT_reg[24]_0 [60]),
        .I3(Q[28]),
        .I4(\CRC_OUT_reg[24]_0 [16]),
        .O(\CRC_OUT[19]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair343" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[19]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [3]),
        .I1(Q[1]),
        .I2(\CRC_OUT_reg[24]_0 [33]),
        .I3(\CRC_OUT_reg[24]_0 [8]),
        .I4(\CRC_OUT[31]_i_4__0_n_0 ),
        .O(\CRC_OUT[19]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair358" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[19]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [47]),
        .I1(Q[15]),
        .I2(\CRC_OUT_reg[24]_0 [29]),
        .O(\CRC_OUT[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[1]_i_1__1 
       (.I0(\CRC_OUT[1]_i_2__0_n_0 ),
        .I1(\CRC_OUT[8]_i_2__0_n_0 ),
        .I2(\CRC_OUT[1]_i_3__0_n_0 ),
        .I3(\CRC_OUT[1]_i_4__0_n_0 ),
        .I4(\CRC_OUT[23]_i_5__0_n_0 ),
        .I5(\CRC_OUT[28]_i_4__0_n_0 ),
        .O(nextCRC32_D64_return056_out));
  (* SOFT_HLUTNM = "soft_lutpair355" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[1]_i_2__0 
       (.I0(\CRC_OUT_reg[24]_0 [62]),
        .I1(Q[30]),
        .I2(\CRC_OUT_reg[24]_0 [49]),
        .I3(Q[17]),
        .O(\CRC_OUT[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[1]_i_3__0 
       (.I0(\CRC_OUT[27]_i_7__0_n_0 ),
        .I1(\CRC_OUT[19]_i_4__0_n_0 ),
        .I2(Q[31]),
        .I3(\CRC_OUT_reg[24]_0 [63]),
        .I4(\CRC_OUT_reg[24]_0 [37]),
        .I5(Q[5]),
        .O(\CRC_OUT[1]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[1]_i_4__0 
       (.I0(\CRC_OUT[23]_i_7__0_n_0 ),
        .I1(\CRC_OUT[17]_i_8__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [9]),
        .I3(\CRC_OUT_reg[24]_0 [28]),
        .I4(\CRC_OUT[25]_i_7__0_n_0 ),
        .I5(\CRC_OUT[18]_i_7__0_n_0 ),
        .O(\CRC_OUT[1]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[20]_i_1__1 
       (.I0(\CRC_OUT[20]_i_2__0_n_0 ),
        .I1(\CRC_OUT[27]_i_3__0_n_0 ),
        .I2(\CRC_OUT[25]_i_5__0_n_0 ),
        .I3(\CRC_OUT[20]_i_3__0_n_0 ),
        .I4(\CRC_OUT[20]_i_4__0_n_0 ),
        .I5(\CRC_OUT[20]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0116_out));
  (* SOFT_HLUTNM = "soft_lutpair368" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[20]_i_2__0 
       (.I0(\CRC_OUT[19]_i_4__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [34]),
        .I2(Q[2]),
        .O(\CRC_OUT[20]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[20]_i_3__0 
       (.I0(\CRC_OUT[4]_i_4__0_n_0 ),
        .I1(\CRC_OUT[0]_i_3__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [17]),
        .I3(\CRC_OUT_reg[24]_0 [25]),
        .I4(\CRC_OUT[23]_i_8__0_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 [9]),
        .O(\CRC_OUT[20]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[20]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [4]),
        .I1(\CRC_OUT_reg[24]_0 [12]),
        .O(\CRC_OUT[20]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[20]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [23]),
        .I1(\CRC_OUT_reg[24]_0 [21]),
        .O(\CRC_OUT[20]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[21]_i_1__1 
       (.I0(\CRC_OUT[28]_i_5__0_n_0 ),
        .I1(\CRC_OUT[30]_i_4__0_n_0 ),
        .I2(\CRC_OUT[21]_i_2__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [24]),
        .I4(\CRC_OUT_reg[24]_0 [26]),
        .I5(\CRC_OUT[21]_i_3__0_n_0 ),
        .O(nextCRC32_D64_return0118_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[21]_i_2__0 
       (.I0(\CRC_OUT[12]_i_5__0_n_0 ),
        .I1(\CRC_OUT[21]_i_4__0_n_0 ),
        .I2(\CRC_OUT[23]_i_3__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [10]),
        .I4(\CRC_OUT_reg[24]_0 [37]),
        .I5(Q[5]),
        .O(\CRC_OUT[21]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair340" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[21]_i_3__0 
       (.I0(\CRC_OUT_reg[24]_0 [13]),
        .I1(\CRC_OUT_reg[24]_0 [5]),
        .O(\CRC_OUT[21]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[21]_i_4__0 
       (.I0(Q[8]),
        .I1(\CRC_OUT_reg[24]_0 [40]),
        .I2(\CRC_OUT_reg[24]_0 [9]),
        .I3(\CRC_OUT_reg[24]_0 [31]),
        .I4(\CRC_OUT_reg[24]_0 [17]),
        .I5(\CRC_OUT_reg[24]_0 [18]),
        .O(\CRC_OUT[21]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[22]_i_1__1 
       (.I0(\CRC_OUT[22]_i_2__0_n_0 ),
        .I1(\CRC_OUT[30]_i_6__0_n_0 ),
        .I2(\CRC_OUT[22]_i_3__0_n_0 ),
        .I3(\CRC_OUT[22]_i_4__0_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [0]),
        .I5(\CRC_OUT[22]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0120_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[22]_i_2__0 
       (.I0(\CRC_OUT[10]_i_4__0_n_0 ),
        .I1(\CRC_OUT[22]_i_6__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [27]),
        .I3(\CRC_OUT_reg[24]_0 [16]),
        .I4(\CRC_OUT[25]_i_7__0_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 [18]),
        .O(\CRC_OUT[22]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[22]_i_3__0 
       (.I0(\CRC_OUT[31]_i_5__0_n_0 ),
        .I1(\CRC_OUT[23]_i_3__0_n_0 ),
        .I2(\CRC_OUT[22]_i_7__0_n_0 ),
        .I3(\CRC_OUT[26]_i_3__0_n_0 ),
        .I4(\CRC_OUT[30]_i_9__0_n_0 ),
        .I5(\CRC_OUT[29]_i_3__0_n_0 ),
        .O(\CRC_OUT[22]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair360" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[22]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [29]),
        .I1(\CRC_OUT_reg[24]_0 [19]),
        .I2(Q[5]),
        .I3(\CRC_OUT_reg[24]_0 [37]),
        .O(\CRC_OUT[22]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair331" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[22]_i_5__0 
       (.I0(Q[4]),
        .I1(\CRC_OUT_reg[24]_0 [36]),
        .I2(\CRC_OUT_reg[24]_0 [9]),
        .I3(\CRC_OUT_reg[24]_0 [31]),
        .I4(\CRC_OUT_reg[24]_0 [14]),
        .O(\CRC_OUT[22]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair361" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[22]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [24]),
        .I1(\CRC_OUT_reg[24]_0 [44]),
        .I2(Q[12]),
        .I3(\CRC_OUT_reg[24]_0 [12]),
        .O(\CRC_OUT[22]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair339" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[22]_i_7__0 
       (.I0(Q[6]),
        .I1(\CRC_OUT_reg[24]_0 [38]),
        .I2(\CRC_OUT_reg[24]_0 [11]),
        .O(\CRC_OUT[22]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[23]_i_1__1 
       (.I0(\CRC_OUT[23]_i_2__1_n_0 ),
        .I1(\CRC_OUT[31]_i_4__0_n_0 ),
        .I2(\CRC_OUT[23]_i_3__0_n_0 ),
        .I3(\CRC_OUT[23]_i_4__0_n_0 ),
        .I4(\CRC_OUT[23]_i_5__0_n_0 ),
        .I5(\CRC_OUT[23]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return0122_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[23]_i_2__1 
       (.I0(\CRC_OUT[29]_i_3__0_n_0 ),
        .I1(\CRC_OUT[19]_i_4__0_n_0 ),
        .I2(\CRC_OUT[23]_i_7__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [20]),
        .I4(\CRC_OUT[23]_i_8__0_n_0 ),
        .I5(\CRC_OUT[26]_i_7__0_n_0 ),
        .O(\CRC_OUT[23]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair368" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[23]_i_3__0 
       (.I0(\CRC_OUT_reg[24]_0 [34]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\CRC_OUT_reg[24]_0 [35]),
        .O(\CRC_OUT[23]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair332" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[23]_i_4__0 
       (.I0(Q[4]),
        .I1(\CRC_OUT_reg[24]_0 [36]),
        .I2(\CRC_OUT_reg[24]_0 [9]),
        .I3(\CRC_OUT_reg[24]_0 [31]),
        .I4(\CRC_OUT[1]_i_2__0_n_0 ),
        .O(\CRC_OUT[23]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[23]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [6]),
        .I1(\CRC_OUT_reg[24]_0 [13]),
        .I2(\CRC_OUT_reg[24]_0 [46]),
        .I3(Q[14]),
        .I4(\CRC_OUT_reg[24]_0 [0]),
        .I5(\CRC_OUT[24]_i_2__1_n_0 ),
        .O(\CRC_OUT[23]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair330" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[23]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [29]),
        .I1(\CRC_OUT_reg[24]_0 [19]),
        .I2(\CRC_OUT_reg[24]_0 [42]),
        .I3(Q[10]),
        .O(\CRC_OUT[23]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[23]_i_7__0 
       (.I0(Q[15]),
        .I1(\CRC_OUT_reg[24]_0 [47]),
        .O(\CRC_OUT[23]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[23]_i_8__0 
       (.I0(Q[7]),
        .I1(\CRC_OUT_reg[24]_0 [39]),
        .O(\CRC_OUT[23]_i_8__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair369" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[24]_i_10__0 
       (.I0(Q[5]),
        .I1(\CRC_OUT_reg[24]_0 [37]),
        .I2(\CRC_OUT_reg[24]_0 [10]),
        .O(\CRC_OUT[24]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair332" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_11__0 
       (.I0(Q[4]),
        .I1(\CRC_OUT_reg[24]_0 [36]),
        .O(\CRC_OUT[24]_i_11__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair353" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_12__0 
       (.I0(\CRC_OUT_reg[24]_0 [43]),
        .I1(Q[11]),
        .O(\CRC_OUT[24]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_1__1 
       (.I0(\CRC_OUT[24]_i_2__1_n_0 ),
        .I1(\CRC_OUT[24]_i_3__1_n_0 ),
        .I2(\CRC_OUT[24]_i_4__1_n_0 ),
        .I3(\CRC_OUT[24]_i_5__0_n_0 ),
        .I4(\CRC_OUT[24]_i_6__0_n_0 ),
        .I5(\CRC_OUT[24]_i_7__0_n_0 ),
        .O(nextCRC32_D64_return0124_out));
  (* SOFT_HLUTNM = "soft_lutpair341" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[24]_i_2__1 
       (.I0(\CRC_OUT_reg[24]_0 [1]),
        .I1(\CRC_OUT_reg[24]_0 [17]),
        .I2(\CRC_OUT_reg[24]_0 [27]),
        .I3(Q[24]),
        .I4(\CRC_OUT_reg[24]_0 [56]),
        .O(\CRC_OUT[24]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_3__1 
       (.I0(Q[8]),
        .I1(\CRC_OUT_reg[24]_0 [40]),
        .I2(Q[31]),
        .I3(\CRC_OUT_reg[24]_0 [63]),
        .I4(\CRC_OUT_reg[24]_0 [28]),
        .I5(\CRC_OUT_reg[24]_0 [30]),
        .O(\CRC_OUT[24]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_4__1 
       (.I0(\CRC_OUT[24]_i_8__0_n_0 ),
        .I1(\CRC_OUT[24]_i_9__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [7]),
        .I3(\CRC_OUT_reg[24]_0 [21]),
        .I4(\CRC_OUT_reg[24]_0 [20]),
        .I5(\CRC_OUT_reg[24]_0 [14]),
        .O(\CRC_OUT[24]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_5__0 
       (.I0(\CRC_OUT[30]_i_9__0_n_0 ),
        .I1(\CRC_OUT[24]_i_10__0_n_0 ),
        .I2(\CRC_OUT[24]_i_11__0_n_0 ),
        .I3(\CRC_OUT[24]_i_12__0_n_0 ),
        .I4(\CRC_OUT[19]_i_4__0_n_0 ),
        .I5(\CRC_OUT[31]_i_11__0_n_0 ),
        .O(\CRC_OUT[24]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair362" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[24]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [2]),
        .I1(\CRC_OUT_reg[24]_0 [18]),
        .I2(\CRC_OUT_reg[24]_0 [39]),
        .I3(Q[7]),
        .O(\CRC_OUT[24]_i_6__0_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[24]_i_7__0 
       (.I0(Q[3]),
        .I1(\CRC_OUT_reg[24]_0 [35]),
        .I2(\CRC_OUT_reg[24]_0 [32]),
        .I3(Q[0]),
        .O(\CRC_OUT[24]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair352" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [51]),
        .I1(Q[19]),
        .O(\CRC_OUT[24]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_9__0 
       (.I0(Q[23]),
        .I1(\CRC_OUT_reg[24]_0 [55]),
        .O(\CRC_OUT[24]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair362" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_10__0 
       (.I0(\CRC_OUT_reg[24]_0 [18]),
        .I1(\CRC_OUT_reg[24]_0 [2]),
        .O(\CRC_OUT[25]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_1__1 
       (.I0(\CRC_OUT[25]_i_2__1_n_0 ),
        .I1(\CRC_OUT[25]_i_3__0_n_0 ),
        .I2(\CRC_OUT[25]_i_4__0_n_0 ),
        .I3(\CRC_OUT[25]_i_5__0_n_0 ),
        .I4(\CRC_OUT[25]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return0126_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[25]_i_2__1 
       (.I0(\CRC_OUT[25]_i_7__0_n_0 ),
        .I1(\CRC_OUT[25]_i_8__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [21]),
        .I3(\CRC_OUT_reg[24]_0 [22]),
        .I4(\CRC_OUT_reg[24]_0 [31]),
        .I5(\CRC_OUT_reg[24]_0 [15]),
        .O(\CRC_OUT[25]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[25]_i_3__0 
       (.I0(\CRC_OUT[22]_i_4__0_n_0 ),
        .I1(\CRC_OUT[25]_i_9__0_n_0 ),
        .I2(\CRC_OUT[30]_i_9__0_n_0 ),
        .I3(\CRC_OUT[11]_i_4__0_n_0 ),
        .I4(\CRC_OUT[25]_i_10__0_n_0 ),
        .I5(\CRC_OUT[1]_i_2__0_n_0 ),
        .O(\CRC_OUT[25]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair339" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [11]),
        .I1(\CRC_OUT_reg[24]_0 [38]),
        .I2(Q[6]),
        .I3(\CRC_OUT_reg[24]_0 [40]),
        .I4(Q[8]),
        .O(\CRC_OUT[25]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair338" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_5__0 
       (.I0(Q[9]),
        .I1(\CRC_OUT_reg[24]_0 [41]),
        .I2(Q[4]),
        .I3(\CRC_OUT_reg[24]_0 [36]),
        .I4(\CRC_OUT[30]_i_11__0_n_0 ),
        .O(\CRC_OUT[25]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair337" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [8]),
        .I1(\CRC_OUT_reg[24]_0 [33]),
        .I2(Q[1]),
        .I3(Q[25]),
        .I4(\CRC_OUT_reg[24]_0 [57]),
        .O(\CRC_OUT[25]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_7__0 
       (.I0(Q[26]),
        .I1(\CRC_OUT_reg[24]_0 [58]),
        .O(\CRC_OUT[25]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [44]),
        .I1(Q[12]),
        .O(\CRC_OUT[25]_i_8__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair341" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[25]_i_9__0 
       (.I0(\CRC_OUT_reg[24]_0 [56]),
        .I1(Q[24]),
        .I2(\CRC_OUT_reg[24]_0 [17]),
        .O(\CRC_OUT[25]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_1__1 
       (.I0(\CRC_OUT[26]_i_2__1_n_0 ),
        .I1(\CRC_OUT[26]_i_3__0_n_0 ),
        .I2(\CRC_OUT[27]_i_3__0_n_0 ),
        .I3(\CRC_OUT[26]_i_4__0_n_0 ),
        .I4(\CRC_OUT[31]_i_5__0_n_0 ),
        .I5(\CRC_OUT[26]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0128_out));
  (* SOFT_HLUTNM = "soft_lutpair365" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[26]_i_2__1 
       (.I0(\CRC_OUT_reg[24]_0 [28]),
        .I1(\CRC_OUT_reg[24]_0 [3]),
        .I2(\CRC_OUT_reg[24]_0 [39]),
        .I3(Q[7]),
        .O(\CRC_OUT[26]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_3__0 
       (.I0(Q[15]),
        .I1(\CRC_OUT_reg[24]_0 [47]),
        .I2(\CRC_OUT_reg[24]_0 [57]),
        .I3(Q[25]),
        .I4(\CRC_OUT_reg[24]_0 [41]),
        .I5(Q[9]),
        .O(\CRC_OUT[26]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_4__0 
       (.I0(\CRC_OUT[26]_i_6__0_n_0 ),
        .I1(\CRC_OUT[28]_i_11__0_n_0 ),
        .I2(\CRC_OUT[1]_i_2__0_n_0 ),
        .I3(\CRC_OUT[26]_i_7__0_n_0 ),
        .I4(\CRC_OUT[5]_i_4__0_n_0 ),
        .I5(\CRC_OUT[26]_i_8__0_n_0 ),
        .O(\CRC_OUT[26]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair335" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[26]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [19]),
        .I1(\CRC_OUT_reg[24]_0 [31]),
        .O(\CRC_OUT[26]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [18]),
        .I1(\CRC_OUT_reg[24]_0 [6]),
        .I2(\CRC_OUT_reg[24]_0 [0]),
        .I3(\CRC_OUT_reg[24]_0 [25]),
        .I4(\CRC_OUT_reg[24]_0 [10]),
        .I5(\CRC_OUT_reg[24]_0 [23]),
        .O(\CRC_OUT[26]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[26]_i_7__0 
       (.I0(\CRC_OUT_reg[24]_0 [38]),
        .I1(Q[6]),
        .O(\CRC_OUT[26]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair346" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[26]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [22]),
        .I1(Q[10]),
        .I2(\CRC_OUT_reg[24]_0 [42]),
        .I3(\CRC_OUT_reg[24]_0 [4]),
        .I4(\CRC_OUT_reg[24]_0 [20]),
        .O(\CRC_OUT[26]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_1__1 
       (.I0(\CRC_OUT[27]_i_2__1_n_0 ),
        .I1(\CRC_OUT[27]_i_3__0_n_0 ),
        .I2(\CRC_OUT[31]_i_8__0_n_0 ),
        .I3(\CRC_OUT[27]_i_4__0_n_0 ),
        .I4(\CRC_OUT[28]_i_5__0_n_0 ),
        .I5(\CRC_OUT[27]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return0130_out));
  (* SOFT_HLUTNM = "soft_lutpair364" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[27]_i_2__1 
       (.I0(\CRC_OUT_reg[24]_0 [21]),
        .I1(\CRC_OUT_reg[24]_0 [5]),
        .I2(\CRC_OUT_reg[24]_0 [4]),
        .I3(\CRC_OUT_reg[24]_0 [20]),
        .O(\CRC_OUT[27]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair366" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[27]_i_3__0 
       (.I0(\CRC_OUT[30]_i_9__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [26]),
        .I2(Q[23]),
        .I3(\CRC_OUT_reg[24]_0 [55]),
        .O(\CRC_OUT[27]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_4__0 
       (.I0(\CRC_OUT[27]_i_6__0_n_0 ),
        .I1(\CRC_OUT[27]_i_7__0_n_0 ),
        .I2(\CRC_OUT[10]_i_3__1_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [1]),
        .I4(\CRC_OUT_reg[24]_0 [24]),
        .I5(\CRC_OUT[27]_i_8__0_n_0 ),
        .O(\CRC_OUT[27]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair330" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[27]_i_5__0 
       (.I0(Q[10]),
        .I1(\CRC_OUT_reg[24]_0 [42]),
        .I2(\CRC_OUT_reg[24]_0 [19]),
        .I3(\CRC_OUT_reg[24]_0 [29]),
        .I4(\CRC_OUT[28]_i_10__0_n_0 ),
        .O(\CRC_OUT[27]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair336" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[27]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [45]),
        .I1(Q[13]),
        .I2(\CRC_OUT_reg[24]_0 [25]),
        .O(\CRC_OUT[27]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair348" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[27]_i_7__0 
       (.I0(Q[21]),
        .I1(\CRC_OUT_reg[24]_0 [53]),
        .I2(\CRC_OUT_reg[24]_0 [7]),
        .O(\CRC_OUT[27]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [39]),
        .I1(Q[7]),
        .I2(Q[18]),
        .I3(\CRC_OUT_reg[24]_0 [50]),
        .I4(\CRC_OUT_reg[24]_0 [60]),
        .I5(Q[28]),
        .O(\CRC_OUT[27]_i_8__0_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_10__0 
       (.I0(\CRC_OUT_reg[24]_0 [63]),
        .I1(Q[31]),
        .I2(\CRC_OUT_reg[24]_0 [40]),
        .I3(Q[8]),
        .O(\CRC_OUT[28]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair345" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_11__0 
       (.I0(\CRC_OUT_reg[24]_0 [54]),
        .I1(Q[22]),
        .I2(\CRC_OUT_reg[24]_0 [59]),
        .I3(Q[27]),
        .O(\CRC_OUT[28]_i_11__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[28]_i_12__0 
       (.I0(Q[17]),
        .I1(\CRC_OUT_reg[24]_0 [49]),
        .O(\CRC_OUT[28]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_1__1 
       (.I0(\CRC_OUT[28]_i_2__1_n_0 ),
        .I1(\CRC_OUT[28]_i_3__0_n_0 ),
        .I2(\CRC_OUT[28]_i_4__0_n_0 ),
        .I3(\CRC_OUT[28]_i_5__0_n_0 ),
        .I4(\CRC_OUT[28]_i_6__0_n_0 ),
        .I5(\CRC_OUT[28]_i_7__0_n_0 ),
        .O(nextCRC32_D64_return0132_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_2__1 
       (.I0(\CRC_OUT[28]_i_8__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [26]),
        .I2(\CRC_OUT_reg[24]_0 [25]),
        .I3(Q[29]),
        .I4(\CRC_OUT_reg[24]_0 [61]),
        .I5(\CRC_OUT[28]_i_9__0_n_0 ),
        .O(\CRC_OUT[28]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_3__0 
       (.I0(\CRC_OUT[28]_i_10__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [6]),
        .I2(\CRC_OUT_reg[24]_0 [2]),
        .I3(\CRC_OUT[28]_i_11__0_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [5]),
        .I5(\CRC_OUT_reg[24]_0 [21]),
        .O(\CRC_OUT[28]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [12]),
        .I1(Q[12]),
        .I2(\CRC_OUT_reg[24]_0 [44]),
        .I3(\CRC_OUT_reg[24]_0 [24]),
        .I4(Q[19]),
        .I5(\CRC_OUT_reg[24]_0 [51]),
        .O(\CRC_OUT[28]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_5__0 
       (.I0(\CRC_OUT[28]_i_12__0_n_0 ),
        .I1(Q[30]),
        .I2(\CRC_OUT_reg[24]_0 [62]),
        .I3(\CRC_OUT_reg[24]_0 [27]),
        .I4(Q[24]),
        .I5(\CRC_OUT_reg[24]_0 [56]),
        .O(\CRC_OUT[28]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair371" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[28]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [20]),
        .I1(\CRC_OUT_reg[24]_0 [22]),
        .O(\CRC_OUT[28]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair344" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[28]_i_7__0 
       (.I0(Q[14]),
        .I1(\CRC_OUT_reg[24]_0 [46]),
        .I2(\CRC_OUT_reg[24]_0 [30]),
        .I3(\CRC_OUT_reg[24]_0 [28]),
        .I4(\CRC_OUT[25]_i_6__0_n_0 ),
        .O(\CRC_OUT[28]_i_7__0_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_8__0 
       (.I0(Q[11]),
        .I1(\CRC_OUT_reg[24]_0 [43]),
        .I2(\CRC_OUT_reg[24]_0 [41]),
        .I3(Q[9]),
        .O(\CRC_OUT[28]_i_8__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair367" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[28]_i_9__0 
       (.I0(Q[18]),
        .I1(\CRC_OUT_reg[24]_0 [50]),
        .O(\CRC_OUT[28]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_1__1 
       (.I0(\CRC_OUT[29]_i_2__1_n_0 ),
        .I1(\CRC_OUT[29]_i_3__0_n_0 ),
        .I2(\CRC_OUT[29]_i_4__0_n_0 ),
        .I3(\CRC_OUT[29]_i_5__0_n_0 ),
        .I4(\CRC_OUT[29]_i_6__0_n_0 ),
        .I5(\CRC_OUT[29]_i_7__0_n_0 ),
        .O(nextCRC32_D64_return0134_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_2__1 
       (.I0(Q[30]),
        .I1(\CRC_OUT_reg[24]_0 [62]),
        .I2(\CRC_OUT[29]_i_8__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [27]),
        .I4(\CRC_OUT_reg[24]_0 [44]),
        .I5(Q[12]),
        .O(\CRC_OUT[29]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair333" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[29]_i_3__0 
       (.I0(\CRC_OUT_reg[24]_0 [55]),
        .I1(Q[23]),
        .I2(\CRC_OUT_reg[24]_0 [26]),
        .O(\CRC_OUT[29]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[29]_i_4__0 
       (.I0(Q[2]),
        .I1(\CRC_OUT_reg[24]_0 [34]),
        .O(\CRC_OUT[29]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [23]),
        .I1(\CRC_OUT_reg[24]_0 [21]),
        .I2(\CRC_OUT[12]_i_2__1_n_0 ),
        .I3(\CRC_OUT[11]_i_4__0_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [6]),
        .I5(\CRC_OUT_reg[24]_0 [13]),
        .O(\CRC_OUT[29]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [29]),
        .I1(\CRC_OUT_reg[24]_0 [22]),
        .I2(Q[10]),
        .I3(\CRC_OUT_reg[24]_0 [42]),
        .I4(\CRC_OUT[30]_i_11__0_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 [7]),
        .O(\CRC_OUT[29]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_7__0 
       (.I0(Q[26]),
        .I1(\CRC_OUT_reg[24]_0 [58]),
        .I2(\CRC_OUT_reg[24]_0 [45]),
        .I3(Q[13]),
        .I4(\CRC_OUT_reg[24]_0 [25]),
        .I5(\CRC_OUT[26]_i_3__0_n_0 ),
        .O(\CRC_OUT[29]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair349" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[29]_i_8__0 
       (.I0(Q[28]),
        .I1(\CRC_OUT_reg[24]_0 [60]),
        .I2(\CRC_OUT_reg[24]_0 [50]),
        .I3(Q[18]),
        .O(\CRC_OUT[29]_i_8__0_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[2]_i_1__1 
       (.I0(\CRC_OUT[2]_i_2__1_n_0 ),
        .I1(\CRC_OUT[11]_i_6__0_n_0 ),
        .I2(\CRC_OUT[2]_i_3__0_n_0 ),
        .O(nextCRC32_D64_return068_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[2]_i_2__1 
       (.I0(\CRC_OUT[30]_i_11__0_n_0 ),
        .I1(\CRC_OUT[5]_i_4__0_n_0 ),
        .I2(\CRC_OUT[15]_i_4__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [16]),
        .I4(\CRC_OUT[2]_i_4__0_n_0 ),
        .I5(\CRC_OUT[26]_i_7__0_n_0 ),
        .O(\CRC_OUT[2]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[2]_i_3__0 
       (.I0(\CRC_OUT[2]_i_5__0_n_0 ),
        .I1(\CRC_OUT[8]_i_5__0_n_0 ),
        .I2(\CRC_OUT[17]_i_6__0_n_0 ),
        .I3(\CRC_OUT[24]_i_6__0_n_0 ),
        .I4(\CRC_OUT[10]_i_3__1_n_0 ),
        .I5(\CRC_OUT[27]_i_7__0_n_0 ),
        .O(\CRC_OUT[2]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair369" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[2]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [37]),
        .I1(Q[5]),
        .O(\CRC_OUT[2]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[2]_i_5__0 
       (.I0(Q[27]),
        .I1(\CRC_OUT_reg[24]_0 [59]),
        .I2(\CRC_OUT_reg[24]_0 [35]),
        .I3(Q[3]),
        .I4(\CRC_OUT_reg[24]_0 [8]),
        .I5(\CRC_OUT_reg[24]_0 [30]),
        .O(\CRC_OUT[2]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair354" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[30]_i_10__0 
       (.I0(Q[31]),
        .I1(\CRC_OUT_reg[24]_0 [63]),
        .O(\CRC_OUT[30]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair352" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[30]_i_11__0 
       (.I0(Q[19]),
        .I1(\CRC_OUT_reg[24]_0 [51]),
        .I2(\CRC_OUT_reg[24]_0 [52]),
        .I3(Q[20]),
        .O(\CRC_OUT[30]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[30]_i_1__1 
       (.I0(\CRC_OUT[30]_i_2__1_n_0 ),
        .I1(\CRC_OUT[30]_i_3__0_n_0 ),
        .I2(\CRC_OUT[30]_i_4__0_n_0 ),
        .I3(\CRC_OUT[30]_i_5__0_n_0 ),
        .I4(\CRC_OUT[30]_i_6__0_n_0 ),
        .I5(\CRC_OUT[30]_i_7__0_n_0 ),
        .O(nextCRC32_D64_return0136_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[30]_i_2__1 
       (.I0(\CRC_OUT[30]_i_8__0_n_0 ),
        .I1(\CRC_OUT[30]_i_9__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [10]),
        .I3(\CRC_OUT_reg[24]_0 [8]),
        .I4(\CRC_OUT[30]_i_10__0_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 [4]),
        .O(\CRC_OUT[30]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[30]_i_3__0 
       (.I0(Q[14]),
        .I1(\CRC_OUT_reg[24]_0 [46]),
        .I2(\CRC_OUT_reg[24]_0 [30]),
        .I3(\CRC_OUT_reg[24]_0 [28]),
        .I4(\CRC_OUT_reg[24]_0 [24]),
        .I5(\CRC_OUT_reg[24]_0 [26]),
        .O(\CRC_OUT[30]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair347" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[30]_i_4__0 
       (.I0(\CRC_OUT[30]_i_11__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [42]),
        .I2(Q[10]),
        .I3(\CRC_OUT_reg[24]_0 [22]),
        .I4(\CRC_OUT_reg[24]_0 [29]),
        .O(\CRC_OUT[30]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair348" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[30]_i_5__0 
       (.I0(\CRC_OUT[10]_i_3__1_n_0 ),
        .I1(Q[21]),
        .I2(\CRC_OUT_reg[24]_0 [53]),
        .I3(\CRC_OUT_reg[24]_0 [7]),
        .I4(\CRC_OUT_reg[24]_0 [14]),
        .O(\CRC_OUT[30]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair342" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[30]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [23]),
        .I1(\CRC_OUT_reg[24]_0 [43]),
        .I2(Q[11]),
        .I3(\CRC_OUT_reg[24]_0 [45]),
        .I4(Q[13]),
        .O(\CRC_OUT[30]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair351" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[30]_i_7__0 
       (.I0(Q[3]),
        .I1(\CRC_OUT_reg[24]_0 [35]),
        .I2(\CRC_OUT_reg[24]_0 [59]),
        .I3(Q[27]),
        .O(\CRC_OUT[30]_i_7__0_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[30]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [56]),
        .I1(Q[24]),
        .I2(\CRC_OUT_reg[24]_0 [27]),
        .O(\CRC_OUT[30]_i_8__0_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[30]_i_9__0 
       (.I0(Q[29]),
        .I1(\CRC_OUT_reg[24]_0 [61]),
        .I2(Q[16]),
        .I3(\CRC_OUT_reg[24]_0 [48]),
        .O(\CRC_OUT[30]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair331" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_10__0 
       (.I0(\CRC_OUT_reg[24]_0 [31]),
        .I1(\CRC_OUT_reg[24]_0 [9]),
        .I2(\CRC_OUT_reg[24]_0 [36]),
        .I3(Q[4]),
        .O(\CRC_OUT[31]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair357" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_11__0 
       (.I0(Q[25]),
        .I1(\CRC_OUT_reg[24]_0 [57]),
        .I2(\CRC_OUT_reg[24]_0 [47]),
        .I3(Q[15]),
        .O(\CRC_OUT[31]_i_11__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair359" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[31]_i_12 
       (.I0(\CRC_OUT_reg[24]_0 [53]),
        .I1(Q[21]),
        .O(\CRC_OUT[31]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \CRC_OUT[31]_i_2__0 
       (.I0(frame_start_del),
        .I1(transmit_pause_frame_valid),
        .O(\CRC_OUT[31]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[31]_i_3__0 
       (.I0(\CRC_OUT[31]_i_4__0_n_0 ),
        .I1(\CRC_OUT[31]_i_5__0_n_0 ),
        .I2(\CRC_OUT[31]_i_6__0_n_0 ),
        .I3(\CRC_OUT[31]_i_7__0_n_0 ),
        .I4(\CRC_OUT[31]_i_8__0_n_0 ),
        .I5(\CRC_OUT[31]_i_9__0_n_0 ),
        .O(nextCRC32_D64_return0138_out));
  (* SOFT_HLUTNM = "soft_lutpair345" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[31]_i_4__0 
       (.I0(Q[27]),
        .I1(\CRC_OUT_reg[24]_0 [59]),
        .I2(Q[22]),
        .I3(\CRC_OUT_reg[24]_0 [54]),
        .I4(\CRC_OUT_reg[24]_0 [15]),
        .O(\CRC_OUT[31]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair356" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_5__0 
       (.I0(Q[28]),
        .I1(\CRC_OUT_reg[24]_0 [60]),
        .I2(\CRC_OUT_reg[24]_0 [52]),
        .I3(Q[20]),
        .O(\CRC_OUT[31]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[31]_i_6__0 
       (.I0(\CRC_OUT[1]_i_2__0_n_0 ),
        .I1(\CRC_OUT[31]_i_10__0_n_0 ),
        .I2(\CRC_OUT[31]_i_11__0_n_0 ),
        .I3(Q[1]),
        .I4(\CRC_OUT_reg[24]_0 [33]),
        .I5(\CRC_OUT_reg[24]_0 [8]),
        .O(\CRC_OUT[31]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[31]_i_7__0 
       (.I0(\CRC_OUT[31]_i_12_n_0 ),
        .I1(\CRC_OUT[5]_i_4__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [29]),
        .I3(\CRC_OUT_reg[24]_0 [25]),
        .I4(\CRC_OUT_reg[24]_0 [27]),
        .I5(\CRC_OUT_reg[24]_0 [5]),
        .O(\CRC_OUT[31]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair353" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_8__0 
       (.I0(\CRC_OUT_reg[24]_0 [23]),
        .I1(\CRC_OUT_reg[24]_0 [43]),
        .I2(Q[11]),
        .I3(\CRC_OUT_reg[24]_0 [11]),
        .O(\CRC_OUT[31]_i_8__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair344" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_9__0 
       (.I0(\CRC_OUT_reg[24]_0 [28]),
        .I1(\CRC_OUT_reg[24]_0 [30]),
        .I2(\CRC_OUT_reg[24]_0 [46]),
        .I3(Q[14]),
        .O(\CRC_OUT[31]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[3]_i_1__1 
       (.I0(\CRC_OUT[7]_i_4__0_n_0 ),
        .I1(\CRC_OUT[3]_i_2__0_n_0 ),
        .I2(\CRC_OUT[3]_i_3__0_n_0 ),
        .I3(\CRC_OUT[24]_i_6__0_n_0 ),
        .I4(\CRC_OUT[19]_i_5__0_n_0 ),
        .I5(\CRC_OUT[31]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return075_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[3]_i_2__0 
       (.I0(Q[8]),
        .I1(\CRC_OUT_reg[24]_0 [40]),
        .I2(\CRC_OUT[27]_i_7__0_n_0 ),
        .I3(\CRC_OUT[10]_i_3__1_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [19]),
        .I5(\CRC_OUT[26]_i_7__0_n_0 ),
        .O(\CRC_OUT[3]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[3]_i_3__0 
       (.I0(\CRC_OUT_reg[24]_0 [14]),
        .I1(\CRC_OUT_reg[24]_0 [31]),
        .I2(\CRC_OUT_reg[24]_0 [9]),
        .I3(\CRC_OUT_reg[24]_0 [36]),
        .I4(Q[4]),
        .I5(\CRC_OUT[24]_i_2__1_n_0 ),
        .O(\CRC_OUT[3]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_1__1 
       (.I0(\CRC_OUT[4]_i_2__1_n_0 ),
        .I1(\CRC_OUT[4]_i_3__0_n_0 ),
        .I2(\CRC_OUT[4]_i_4__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [3]),
        .I4(\CRC_OUT[29]_i_7__0_n_0 ),
        .I5(\CRC_OUT[18]_i_5__0_n_0 ),
        .O(nextCRC32_D64_return080_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_2__1 
       (.I0(\CRC_OUT[18]_i_7__0_n_0 ),
        .I1(\CRC_OUT[14]_i_5__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [31]),
        .I3(\CRC_OUT_reg[24]_0 [15]),
        .I4(\CRC_OUT_reg[24]_0 [30]),
        .I5(\CRC_OUT_reg[24]_0 [6]),
        .O(\CRC_OUT[4]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_3__0 
       (.I0(\CRC_OUT[28]_i_10__0_n_0 ),
        .I1(\CRC_OUT[24]_i_6__0_n_0 ),
        .I2(\CRC_OUT[11]_i_3__0_n_0 ),
        .I3(\CRC_OUT[22]_i_6__0_n_0 ),
        .I4(\CRC_OUT[16]_i_5__0_n_0 ),
        .I5(\CRC_OUT[22]_i_7__0_n_0 ),
        .O(\CRC_OUT[4]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair337" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[4]_i_4__0 
       (.I0(Q[1]),
        .I1(\CRC_OUT_reg[24]_0 [33]),
        .I2(\CRC_OUT_reg[24]_0 [8]),
        .O(\CRC_OUT[4]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[5]_i_1__1 
       (.I0(\CRC_OUT[5]_i_2__1_n_0 ),
        .I1(\CRC_OUT[5]_i_3__0_n_0 ),
        .I2(\CRC_OUT[5]_i_4__0_n_0 ),
        .I3(\CRC_OUT[5]_i_5__0_n_0 ),
        .I4(\CRC_OUT[27]_i_5__0_n_0 ),
        .I5(\CRC_OUT[5]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return086_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[5]_i_2__1 
       (.I0(\CRC_OUT[26]_i_2__1_n_0 ),
        .I1(\CRC_OUT[13]_i_4__0_n_0 ),
        .I2(\CRC_OUT[27]_i_7__0_n_0 ),
        .I3(\CRC_OUT[28]_i_11__0_n_0 ),
        .I4(\CRC_OUT[27]_i_2__1_n_0 ),
        .I5(\CRC_OUT[24]_i_10__0_n_0 ),
        .O(\CRC_OUT[5]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair338" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[5]_i_3__0 
       (.I0(Q[9]),
        .I1(\CRC_OUT_reg[24]_0 [41]),
        .O(\CRC_OUT[5]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair361" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[5]_i_4__0 
       (.I0(Q[12]),
        .I1(\CRC_OUT_reg[24]_0 [44]),
        .I2(\CRC_OUT_reg[24]_0 [24]),
        .O(\CRC_OUT[5]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[5]_i_5__0 
       (.I0(\CRC_OUT[28]_i_12__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [61]),
        .I2(Q[29]),
        .I3(\CRC_OUT[28]_i_9__0_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [51]),
        .I5(Q[19]),
        .O(\CRC_OUT[5]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair334" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[5]_i_6__0 
       (.I0(\CRC_OUT_reg[24]_0 [0]),
        .I1(Q[14]),
        .I2(\CRC_OUT_reg[24]_0 [46]),
        .I3(\CRC_OUT_reg[24]_0 [13]),
        .I4(\CRC_OUT_reg[24]_0 [6]),
        .O(\CRC_OUT[5]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[6]_i_1__1 
       (.I0(\CRC_OUT[6]_i_2__1_n_0 ),
        .I1(\CRC_OUT[6]_i_3__0_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [30]),
        .I3(\CRC_OUT_reg[24]_0 [8]),
        .I4(\CRC_OUT[29]_i_6__0_n_0 ),
        .I5(\CRC_OUT[25]_i_4__0_n_0 ),
        .O(nextCRC32_D64_return091_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[6]_i_2__1 
       (.I0(Q[30]),
        .I1(\CRC_OUT_reg[24]_0 [62]),
        .I2(\CRC_OUT[29]_i_8__0_n_0 ),
        .I3(\CRC_OUT[23]_i_7__0_n_0 ),
        .I4(\CRC_OUT_reg[24]_0 [14]),
        .I5(\CRC_OUT[7]_i_5__0_n_0 ),
        .O(\CRC_OUT[6]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[6]_i_3__0 
       (.I0(\CRC_OUT[27]_i_2__1_n_0 ),
        .I1(\CRC_OUT[13]_i_4__0_n_0 ),
        .I2(\CRC_OUT[28]_i_8__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [2]),
        .I4(\CRC_OUT_reg[24]_0 [6]),
        .I5(\CRC_OUT[27]_i_6__0_n_0 ),
        .O(\CRC_OUT[6]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[7]_i_1__1 
       (.I0(\CRC_OUT[7]_i_2__1_n_0 ),
        .I1(\CRC_OUT[7]_i_3__0_n_0 ),
        .I2(\CRC_OUT[20]_i_2__0_n_0 ),
        .I3(\CRC_OUT[29]_i_6__0_n_0 ),
        .I4(\CRC_OUT[7]_i_4__0_n_0 ),
        .O(nextCRC32_D64_return093_out));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[7]_i_2__1 
       (.I0(\CRC_OUT[7]_i_5__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [8]),
        .I2(\CRC_OUT_reg[24]_0 [2]),
        .I3(\CRC_OUT_reg[24]_0 [24]),
        .I4(\CRC_OUT_reg[24]_0 [15]),
        .O(\CRC_OUT[7]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[7]_i_3__0 
       (.I0(\CRC_OUT[26]_i_3__0_n_0 ),
        .I1(\CRC_OUT[26]_i_2__1_n_0 ),
        .I2(\CRC_OUT[16]_i_4__1_n_0 ),
        .I3(\CRC_OUT[10]_i_3__1_n_0 ),
        .I4(\CRC_OUT[16]_i_5__0_n_0 ),
        .I5(\CRC_OUT[9]_i_6__0_n_0 ),
        .O(\CRC_OUT[7]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[7]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [10]),
        .I1(\CRC_OUT_reg[24]_0 [37]),
        .I2(Q[5]),
        .I3(\CRC_OUT_reg[24]_0 [25]),
        .I4(Q[13]),
        .I5(\CRC_OUT_reg[24]_0 [45]),
        .O(\CRC_OUT[7]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair350" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[7]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [54]),
        .I1(Q[22]),
        .I2(\CRC_OUT_reg[24]_0 [56]),
        .I3(Q[24]),
        .O(\CRC_OUT[7]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_1__1 
       (.I0(\CRC_OUT[8]_i_2__0_n_0 ),
        .I1(\CRC_OUT[20]_i_4__0_n_0 ),
        .I2(\CRC_OUT[8]_i_3__0_n_0 ),
        .I3(\CRC_OUT[8]_i_4__0_n_0 ),
        .I4(\CRC_OUT[25]_i_6__0_n_0 ),
        .I5(\CRC_OUT[30]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return094_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_2__0 
       (.I0(\CRC_OUT_reg[24]_0 [35]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(\CRC_OUT_reg[24]_0 [34]),
        .I4(\CRC_OUT_reg[24]_0 [11]),
        .I5(\CRC_OUT[26]_i_7__0_n_0 ),
        .O(\CRC_OUT[8]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_3__0 
       (.I0(\CRC_OUT[28]_i_10__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [22]),
        .I2(\CRC_OUT[12]_i_6__0_n_0 ),
        .I3(\CRC_OUT[30]_i_11__0_n_0 ),
        .I4(\CRC_OUT[24]_i_10__0_n_0 ),
        .I5(\CRC_OUT[16]_i_5__0_n_0 ),
        .O(\CRC_OUT[8]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_4__0 
       (.I0(\CRC_OUT[11]_i_4__0_n_0 ),
        .I1(\CRC_OUT[8]_i_5__0_n_0 ),
        .I2(\CRC_OUT[8]_i_6__0_n_0 ),
        .I3(\CRC_OUT_reg[24]_0 [31]),
        .I4(\CRC_OUT[28]_i_11__0_n_0 ),
        .I5(\CRC_OUT[29]_i_8__0_n_0 ),
        .O(\CRC_OUT[8]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[8]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [17]),
        .I1(\CRC_OUT_reg[24]_0 [1]),
        .O(\CRC_OUT[8]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair363" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[8]_i_6__0 
       (.I0(Q[0]),
        .I1(\CRC_OUT_reg[24]_0 [32]),
        .O(\CRC_OUT[8]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_1__1 
       (.I0(\CRC_OUT[9]_i_2__1_n_0 ),
        .I1(\CRC_OUT[9]_i_3__0_n_0 ),
        .I2(\CRC_OUT[9]_i_4__0_n_0 ),
        .I3(\CRC_OUT[12]_i_5__0_n_0 ),
        .I4(\CRC_OUT[25]_i_5__0_n_0 ),
        .I5(\CRC_OUT[19]_i_6__0_n_0 ),
        .O(nextCRC32_D64_return096_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_2__1 
       (.I0(\CRC_OUT[18]_i_6__0_n_0 ),
        .I1(\CRC_OUT[10]_i_3__1_n_0 ),
        .I2(\CRC_OUT_reg[24]_0 [9]),
        .I3(\CRC_OUT_reg[24]_0 [4]),
        .I4(\CRC_OUT[17]_i_8__0_n_0 ),
        .I5(\CRC_OUT[9]_i_5__0_n_0 ),
        .O(\CRC_OUT[9]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_3__0 
       (.I0(\CRC_OUT[24]_i_6__0_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 [55]),
        .I2(Q[23]),
        .I3(\CRC_OUT_reg[24]_0 [1]),
        .I4(\CRC_OUT[22]_i_6__0_n_0 ),
        .I5(\CRC_OUT[9]_i_6__0_n_0 ),
        .O(\CRC_OUT[9]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_4__0 
       (.I0(\CRC_OUT_reg[24]_0 [5]),
        .I1(\CRC_OUT_reg[24]_0 [13]),
        .I2(Q[6]),
        .I3(\CRC_OUT_reg[24]_0 [38]),
        .I4(\CRC_OUT_reg[24]_0 [11]),
        .I5(\CRC_OUT[23]_i_3__0_n_0 ),
        .O(\CRC_OUT[9]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair356" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[9]_i_5__0 
       (.I0(\CRC_OUT_reg[24]_0 [60]),
        .I1(Q[28]),
        .O(\CRC_OUT[9]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair342" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[9]_i_6__0 
       (.I0(Q[11]),
        .I1(\CRC_OUT_reg[24]_0 [43]),
        .I2(\CRC_OUT_reg[24]_0 [23]),
        .O(\CRC_OUT[9]_i_6__0_n_0 ));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[0] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0),
        .Q(Q[0]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[10] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return098_out),
        .Q(Q[10]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[11] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0100_out),
        .Q(Q[11]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[12] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0102_out),
        .Q(Q[12]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[13] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0104_out),
        .Q(Q[13]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[14] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0106_out),
        .Q(Q[14]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[15] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0108_out),
        .Q(Q[15]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[16] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0109_out),
        .Q(Q[16]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[17] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0110_out),
        .Q(Q[17]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[18] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0112_out),
        .Q(Q[18]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[19] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0114_out),
        .Q(Q[19]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[1] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return056_out),
        .Q(Q[1]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[20] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0116_out),
        .Q(Q[20]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[21] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0118_out),
        .Q(Q[21]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[22] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0120_out),
        .Q(Q[22]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[23] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0122_out),
        .Q(Q[23]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[24] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0124_out),
        .Q(Q[24]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[25] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0126_out),
        .Q(Q[25]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[26] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0128_out),
        .Q(Q[26]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[27] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0130_out),
        .Q(Q[27]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[28] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0132_out),
        .Q(Q[28]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[29] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0134_out),
        .Q(Q[29]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[2] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return068_out),
        .Q(Q[2]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[30] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0136_out),
        .Q(Q[30]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[31] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return0138_out),
        .Q(Q[31]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[3] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return075_out),
        .Q(Q[3]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[4] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return080_out),
        .Q(Q[4]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[5] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return086_out),
        .Q(Q[5]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[6] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return091_out),
        .Q(Q[6]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[7] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return093_out),
        .Q(Q[7]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[8] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return094_out),
        .Q(Q[8]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[9] 
       (.C(clk_i),
        .CE(\CRC_OUT[31]_i_2__0_n_0 ),
        .D(nextCRC32_D64_return096_out),
        .Q(Q[9]),
        .S(SS));
endmodule

(* ORIG_REF_NAME = "CRC32_D64" *) 
module switch_elements_CRC32_D64_3
   (\CRC_OUT_reg[29]_0 ,
    \CRC_OUT_reg[29]_1 ,
    \CRC_OUT_reg[25]_0 ,
    \rxd64_d3_reg[37] ,
    \CRC_OUT_reg[11]_0 ,
    Q,
    \CRC_OUT_reg[18]_0 ,
    \rxd64_d3_reg[48] ,
    \CRC_OUT_reg[14]_0 ,
    \CRC_OUT_reg[7]_0 ,
    \CRC_OUT_reg[17]_0 ,
    \CRC_OUT_reg[27]_0 ,
    \rxd64_d3_reg[54] ,
    \CRC_OUT_reg[15]_0 ,
    \CRC_OUT_reg[26]_0 ,
    \CRC_OUT_reg[30]_0 ,
    \CRC_OUT_reg[28]_0 ,
    \CRC_OUT_reg[15]_1 ,
    \CRC_OUT_reg[28]_1 ,
    \CRC_OUT_reg[28]_2 ,
    \CRC_OUT_reg[15]_2 ,
    \CRC_OUT_reg[2]_0 ,
    \CRC_OUT_reg[26]_1 ,
    \rxd64_d3_reg[2] ,
    \rxd64_d3_reg[33] ,
    \CRC_OUT_reg[10]_0 ,
    \CRC_OUT_reg[19]_0 ,
    \CRC_OUT_reg[30]_1 ,
    \CRC_OUT_reg[30]_2 ,
    \CRC_OUT_reg[9]_0 ,
    \CRC_OUT_reg[3]_0 ,
    \CRC_OUT_reg[22]_0 ,
    \CRC_OUT_reg[20]_0 ,
    \CRC_OUT_reg[29]_2 ,
    \CRC_OUT_reg[3]_1 ,
    \CRC_OUT_reg[0]_0 ,
    \CRC_OUT_reg[31]_0 ,
    \CRC_OUT_reg[16]_0 ,
    \rxd64_d3_reg[37]_0 ,
    \CRC_OUT_reg[9]_1 ,
    \CRC_OUT_reg[23]_0 ,
    \CRC_OUT_reg[24]_0 ,
    \CRC_OUT_reg[24]_1 ,
    \CRC_OUT_reg[24]_2 ,
    rxd64_d3,
    \CRC_OUT_reg[1]_0 ,
    \CRC_OUT_reg[6]_0 ,
    \CRC_OUT_reg[22]_1 ,
    \CRC_OUT_reg[22]_2 ,
    \CRC_OUT_reg[29]_3 ,
    \CRC_OUT_reg[29]_4 ,
    \CRC_OUT_reg[29]_5 ,
    SS,
    E,
    \CRC_OUT_reg[31]_1 ,
    clk_i);
  output \CRC_OUT_reg[29]_0 ;
  output \CRC_OUT_reg[29]_1 ;
  output \CRC_OUT_reg[25]_0 ;
  output \rxd64_d3_reg[37] ;
  output \CRC_OUT_reg[11]_0 ;
  output [31:0]Q;
  output \CRC_OUT_reg[18]_0 ;
  output \rxd64_d3_reg[48] ;
  output \CRC_OUT_reg[14]_0 ;
  output \CRC_OUT_reg[7]_0 ;
  output \CRC_OUT_reg[17]_0 ;
  output \CRC_OUT_reg[27]_0 ;
  output \rxd64_d3_reg[54] ;
  output \CRC_OUT_reg[15]_0 ;
  output \CRC_OUT_reg[26]_0 ;
  output \CRC_OUT_reg[30]_0 ;
  output \CRC_OUT_reg[28]_0 ;
  output \CRC_OUT_reg[15]_1 ;
  output \CRC_OUT_reg[28]_1 ;
  output \CRC_OUT_reg[28]_2 ;
  output \CRC_OUT_reg[15]_2 ;
  output \CRC_OUT_reg[2]_0 ;
  output \CRC_OUT_reg[26]_1 ;
  output \rxd64_d3_reg[2] ;
  output \rxd64_d3_reg[33] ;
  output \CRC_OUT_reg[10]_0 ;
  output \CRC_OUT_reg[19]_0 ;
  output \CRC_OUT_reg[30]_1 ;
  output \CRC_OUT_reg[30]_2 ;
  output \CRC_OUT_reg[9]_0 ;
  output \CRC_OUT_reg[3]_0 ;
  output \CRC_OUT_reg[22]_0 ;
  output \CRC_OUT_reg[20]_0 ;
  output \CRC_OUT_reg[29]_2 ;
  output \CRC_OUT_reg[3]_1 ;
  output \CRC_OUT_reg[0]_0 ;
  output \CRC_OUT_reg[31]_0 ;
  output \CRC_OUT_reg[16]_0 ;
  output \rxd64_d3_reg[37]_0 ;
  output \CRC_OUT_reg[9]_1 ;
  output \CRC_OUT_reg[23]_0 ;
  input \CRC_OUT_reg[24]_0 ;
  input \CRC_OUT_reg[24]_1 ;
  input \CRC_OUT_reg[24]_2 ;
  input [36:0]rxd64_d3;
  input \CRC_OUT_reg[1]_0 ;
  input \CRC_OUT_reg[6]_0 ;
  input \CRC_OUT_reg[22]_1 ;
  input \CRC_OUT_reg[22]_2 ;
  input \CRC_OUT_reg[29]_3 ;
  input \CRC_OUT_reg[29]_4 ;
  input \CRC_OUT_reg[29]_5 ;
  input [0:0]SS;
  input [0:0]E;
  input [30:0]\CRC_OUT_reg[31]_1 ;
  input clk_i;

  wire \CRC_OUT[24]_i_11_n_0 ;
  wire \CRC_OUT[29]_i_2_n_0 ;
  wire \CRC_OUT_reg[0]_0 ;
  wire \CRC_OUT_reg[10]_0 ;
  wire \CRC_OUT_reg[11]_0 ;
  wire \CRC_OUT_reg[14]_0 ;
  wire \CRC_OUT_reg[15]_0 ;
  wire \CRC_OUT_reg[15]_1 ;
  wire \CRC_OUT_reg[15]_2 ;
  wire \CRC_OUT_reg[16]_0 ;
  wire \CRC_OUT_reg[17]_0 ;
  wire \CRC_OUT_reg[18]_0 ;
  wire \CRC_OUT_reg[19]_0 ;
  wire \CRC_OUT_reg[1]_0 ;
  wire \CRC_OUT_reg[20]_0 ;
  wire \CRC_OUT_reg[22]_0 ;
  wire \CRC_OUT_reg[22]_1 ;
  wire \CRC_OUT_reg[22]_2 ;
  wire \CRC_OUT_reg[23]_0 ;
  wire \CRC_OUT_reg[24]_0 ;
  wire \CRC_OUT_reg[24]_1 ;
  wire \CRC_OUT_reg[24]_2 ;
  wire \CRC_OUT_reg[25]_0 ;
  wire \CRC_OUT_reg[26]_0 ;
  wire \CRC_OUT_reg[26]_1 ;
  wire \CRC_OUT_reg[27]_0 ;
  wire \CRC_OUT_reg[28]_0 ;
  wire \CRC_OUT_reg[28]_1 ;
  wire \CRC_OUT_reg[28]_2 ;
  wire \CRC_OUT_reg[29]_0 ;
  wire \CRC_OUT_reg[29]_1 ;
  wire \CRC_OUT_reg[29]_2 ;
  wire \CRC_OUT_reg[29]_3 ;
  wire \CRC_OUT_reg[29]_4 ;
  wire \CRC_OUT_reg[29]_5 ;
  wire \CRC_OUT_reg[2]_0 ;
  wire \CRC_OUT_reg[30]_0 ;
  wire \CRC_OUT_reg[30]_1 ;
  wire \CRC_OUT_reg[30]_2 ;
  wire \CRC_OUT_reg[31]_0 ;
  wire [30:0]\CRC_OUT_reg[31]_1 ;
  wire \CRC_OUT_reg[3]_0 ;
  wire \CRC_OUT_reg[3]_1 ;
  wire \CRC_OUT_reg[6]_0 ;
  wire \CRC_OUT_reg[7]_0 ;
  wire \CRC_OUT_reg[9]_0 ;
  wire \CRC_OUT_reg[9]_1 ;
  wire [0:0]E;
  wire [31:0]Q;
  wire [0:0]SS;
  wire clk_i;
  wire nextCRC32_D64_return0134_out;
  wire [36:0]rxd64_d3;
  wire \rxd64_d3_reg[2] ;
  wire \rxd64_d3_reg[33] ;
  wire \rxd64_d3_reg[37] ;
  wire \rxd64_d3_reg[37]_0 ;
  wire \rxd64_d3_reg[48] ;
  wire \rxd64_d3_reg[54] ;

  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[10]_i_4 
       (.I0(Q[30]),
        .I1(rxd64_d3[1]),
        .O(\CRC_OUT_reg[30]_2 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[12]_i_4 
       (.I0(\CRC_OUT_reg[10]_0 ),
        .I1(\CRC_OUT_reg[19]_0 ),
        .I2(rxd64_d3[28]),
        .I3(rxd64_d3[33]),
        .I4(\CRC_OUT_reg[17]_0 ),
        .I5(\CRC_OUT_reg[18]_0 ),
        .O(\rxd64_d3_reg[33] ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[12]_i_5 
       (.I0(Q[29]),
        .I1(rxd64_d3[2]),
        .I2(Q[21]),
        .I3(rxd64_d3[10]),
        .O(\CRC_OUT_reg[29]_2 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[12]_i_6 
       (.I0(Q[10]),
        .I1(rxd64_d3[21]),
        .O(\CRC_OUT_reg[10]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[13]_i_7 
       (.I0(Q[22]),
        .I1(rxd64_d3[9]),
        .O(\CRC_OUT_reg[22]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_5 
       (.I0(Q[15]),
        .I1(rxd64_d3[16]),
        .I2(rxd64_d3[6]),
        .I3(Q[25]),
        .I4(Q[16]),
        .I5(rxd64_d3[15]),
        .O(\CRC_OUT_reg[15]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_7 
       (.I0(Q[20]),
        .I1(rxd64_d3[11]),
        .O(\CRC_OUT_reg[20]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[18]_i_4 
       (.I0(\CRC_OUT_reg[14]_0 ),
        .I1(\CRC_OUT_reg[7]_0 ),
        .I2(rxd64_d3[34]),
        .I3(rxd64_d3[29]),
        .I4(\CRC_OUT_reg[17]_0 ),
        .I5(\CRC_OUT_reg[27]_0 ),
        .O(\rxd64_d3_reg[48] ));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[18]_i_5 
       (.I0(Q[16]),
        .I1(rxd64_d3[15]),
        .I2(rxd64_d3[13]),
        .I3(Q[18]),
        .O(\CRC_OUT_reg[16]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_6 
       (.I0(Q[14]),
        .I1(rxd64_d3[17]),
        .O(\CRC_OUT_reg[14]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_7 
       (.I0(Q[27]),
        .I1(rxd64_d3[4]),
        .O(\CRC_OUT_reg[27]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[1]_i_4 
       (.I0(\CRC_OUT_reg[15]_0 ),
        .I1(\CRC_OUT_reg[1]_0 ),
        .I2(rxd64_d3[36]),
        .I3(rxd64_d3[29]),
        .I4(\CRC_OUT_reg[26]_0 ),
        .I5(\CRC_OUT_reg[27]_0 ),
        .O(\rxd64_d3_reg[54] ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[22]_i_3 
       (.I0(\CRC_OUT_reg[28]_2 ),
        .I1(\CRC_OUT_reg[22]_1 ),
        .I2(\CRC_OUT_reg[22]_2 ),
        .I3(\CRC_OUT_reg[15]_2 ),
        .I4(\CRC_OUT_reg[29]_1 ),
        .I5(\CRC_OUT_reg[29]_3 ),
        .O(\CRC_OUT_reg[28]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[23]_i_7 
       (.I0(Q[15]),
        .I1(rxd64_d3[16]),
        .O(\CRC_OUT_reg[15]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[23]_i_8 
       (.I0(Q[7]),
        .I1(rxd64_d3[23]),
        .O(\CRC_OUT_reg[7]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_11 
       (.I0(Q[4]),
        .I1(rxd64_d3[24]),
        .O(\CRC_OUT[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_5 
       (.I0(\CRC_OUT_reg[29]_1 ),
        .I1(\CRC_OUT_reg[24]_0 ),
        .I2(\CRC_OUT[24]_i_11_n_0 ),
        .I3(\CRC_OUT_reg[24]_1 ),
        .I4(\CRC_OUT_reg[24]_2 ),
        .I5(\CRC_OUT_reg[25]_0 ),
        .O(\CRC_OUT_reg[29]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[24]_i_7 
       (.I0(Q[3]),
        .I1(rxd64_d3[25]),
        .I2(rxd64_d3[27]),
        .I3(Q[0]),
        .O(\CRC_OUT_reg[3]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_9 
       (.I0(Q[23]),
        .I1(rxd64_d3[8]),
        .O(\CRC_OUT_reg[23]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_5 
       (.I0(Q[9]),
        .I1(rxd64_d3[22]),
        .I2(Q[4]),
        .I3(rxd64_d3[24]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .O(\CRC_OUT_reg[9]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_7 
       (.I0(Q[26]),
        .I1(rxd64_d3[5]),
        .O(\CRC_OUT_reg[26]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_3 
       (.I0(Q[15]),
        .I1(rxd64_d3[16]),
        .I2(rxd64_d3[6]),
        .I3(Q[25]),
        .I4(rxd64_d3[22]),
        .I5(Q[9]),
        .O(\CRC_OUT_reg[15]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[27]_i_3 
       (.I0(\CRC_OUT_reg[29]_1 ),
        .I1(rxd64_d3[31]),
        .I2(Q[23]),
        .I3(rxd64_d3[8]),
        .O(\rxd64_d3_reg[37]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[28]_i_12 
       (.I0(Q[17]),
        .I1(rxd64_d3[14]),
        .O(\CRC_OUT_reg[17]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_2 
       (.I0(\CRC_OUT_reg[11]_0 ),
        .I1(rxd64_d3[31]),
        .I2(rxd64_d3[32]),
        .I3(Q[29]),
        .I4(rxd64_d3[2]),
        .I5(\CRC_OUT_reg[18]_0 ),
        .O(\rxd64_d3_reg[37] ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_5 
       (.I0(\CRC_OUT_reg[17]_0 ),
        .I1(Q[30]),
        .I2(rxd64_d3[1]),
        .I3(rxd64_d3[30]),
        .I4(Q[24]),
        .I5(rxd64_d3[7]),
        .O(\CRC_OUT_reg[30]_1 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_8 
       (.I0(Q[11]),
        .I1(rxd64_d3[20]),
        .I2(rxd64_d3[22]),
        .I3(Q[9]),
        .O(\CRC_OUT_reg[11]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[28]_i_9 
       (.I0(Q[18]),
        .I1(rxd64_d3[13]),
        .O(\CRC_OUT_reg[18]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_1 
       (.I0(\CRC_OUT[29]_i_2_n_0 ),
        .I1(\CRC_OUT_reg[29]_3 ),
        .I2(\CRC_OUT_reg[2]_0 ),
        .I3(\CRC_OUT_reg[29]_4 ),
        .I4(\CRC_OUT_reg[29]_5 ),
        .I5(\CRC_OUT_reg[26]_1 ),
        .O(nextCRC32_D64_return0134_out));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_2 
       (.I0(Q[30]),
        .I1(rxd64_d3[1]),
        .I2(\CRC_OUT_reg[28]_0 ),
        .I3(rxd64_d3[30]),
        .I4(rxd64_d3[19]),
        .I5(Q[12]),
        .O(\CRC_OUT[29]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[29]_i_4 
       (.I0(Q[2]),
        .I1(rxd64_d3[26]),
        .O(\CRC_OUT_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_7 
       (.I0(Q[26]),
        .I1(rxd64_d3[5]),
        .I2(rxd64_d3[18]),
        .I3(Q[13]),
        .I4(rxd64_d3[32]),
        .I5(\CRC_OUT_reg[15]_2 ),
        .O(\CRC_OUT_reg[26]_1 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[29]_i_8 
       (.I0(Q[28]),
        .I1(rxd64_d3[3]),
        .I2(rxd64_d3[13]),
        .I3(Q[18]),
        .O(\CRC_OUT_reg[28]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[30]_i_10 
       (.I0(Q[31]),
        .I1(rxd64_d3[0]),
        .O(\CRC_OUT_reg[31]_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[30]_i_11 
       (.I0(Q[19]),
        .I1(rxd64_d3[12]),
        .I2(rxd64_d3[11]),
        .I3(Q[20]),
        .O(\CRC_OUT_reg[19]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[30]_i_7 
       (.I0(Q[3]),
        .I1(rxd64_d3[25]),
        .I2(rxd64_d3[4]),
        .I3(Q[27]),
        .O(\CRC_OUT_reg[3]_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[30]_i_9 
       (.I0(Q[29]),
        .I1(rxd64_d3[2]),
        .I2(Q[16]),
        .I3(rxd64_d3[15]),
        .O(\CRC_OUT_reg[29]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_10 
       (.I0(Q[25]),
        .I1(rxd64_d3[6]),
        .I2(rxd64_d3[16]),
        .I3(Q[15]),
        .O(\CRC_OUT_reg[25]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_4 
       (.I0(Q[28]),
        .I1(rxd64_d3[3]),
        .I2(rxd64_d3[11]),
        .I3(Q[20]),
        .O(\CRC_OUT_reg[28]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[5]_i_3 
       (.I0(Q[9]),
        .I1(rxd64_d3[22]),
        .O(\CRC_OUT_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[5]_i_5 
       (.I0(\CRC_OUT_reg[17]_0 ),
        .I1(rxd64_d3[2]),
        .I2(Q[29]),
        .I3(\CRC_OUT_reg[18]_0 ),
        .I4(rxd64_d3[12]),
        .I5(Q[19]),
        .O(\rxd64_d3_reg[2] ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[6]_i_2 
       (.I0(Q[30]),
        .I1(rxd64_d3[1]),
        .I2(\CRC_OUT_reg[28]_0 ),
        .I3(\CRC_OUT_reg[15]_0 ),
        .I4(rxd64_d3[35]),
        .I5(\CRC_OUT_reg[6]_0 ),
        .O(\CRC_OUT_reg[30]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[8]_i_6 
       (.I0(Q[0]),
        .I1(rxd64_d3[27]),
        .O(\CRC_OUT_reg[0]_0 ));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[0] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [0]),
        .Q(Q[0]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[10] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [10]),
        .Q(Q[10]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[11] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [11]),
        .Q(Q[11]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[12] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [12]),
        .Q(Q[12]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[13] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [13]),
        .Q(Q[13]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[14] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [14]),
        .Q(Q[14]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[15] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [15]),
        .Q(Q[15]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[16] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [16]),
        .Q(Q[16]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[17] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [17]),
        .Q(Q[17]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[18] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [18]),
        .Q(Q[18]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[19] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [19]),
        .Q(Q[19]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[1] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [1]),
        .Q(Q[1]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[20] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [20]),
        .Q(Q[20]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[21] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [21]),
        .Q(Q[21]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[22] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [22]),
        .Q(Q[22]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[23] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [23]),
        .Q(Q[23]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[24] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [24]),
        .Q(Q[24]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[25] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [25]),
        .Q(Q[25]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[26] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [26]),
        .Q(Q[26]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[27] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [27]),
        .Q(Q[27]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[28] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [28]),
        .Q(Q[28]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[29] 
       (.C(clk_i),
        .CE(E),
        .D(nextCRC32_D64_return0134_out),
        .Q(Q[29]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[2] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [2]),
        .Q(Q[2]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[30] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [29]),
        .Q(Q[30]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[31] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [30]),
        .Q(Q[31]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[3] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [3]),
        .Q(Q[3]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[4] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [4]),
        .Q(Q[4]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[5] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [5]),
        .Q(Q[5]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[6] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [6]),
        .Q(Q[6]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[7] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [7]),
        .Q(Q[7]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[8] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [8]),
        .Q(Q[8]),
        .S(SS));
  FDSE #(
    .INIT(1'b1)) 
    \CRC_OUT_reg[9] 
       (.C(clk_i),
        .CE(E),
        .D(\CRC_OUT_reg[31]_1 [9]),
        .Q(Q[9]),
        .S(SS));
endmodule

(* ORIG_REF_NAME = "CRC32_D8" *) 
module switch_elements_CRC32_D8
   (D,
    E,
    \TX_DATA_VALID_DEL13_reg[7] ,
    \TX_DATA_DEL14_reg[32] ,
    fcs_enabled_int,
    TX_DATA_VALID_DEL13,
    \TX_DATA_DEL14_reg[58] ,
    TX_DATA_DEL13,
    \TX_DATA_DEL14_reg[50] ,
    \TX_DATA_DEL14_reg[33] ,
    \TX_DATA_DEL14_reg[26] ,
    \OVERFLOW_DATA_reg[8] ,
    \TX_DATA_DEL14_reg[21] ,
    Q,
    \OVERFLOW_DATA_reg[2] ,
    txstatplus_int,
    \OVERFLOW_DATA_reg[2]_0 ,
    TX_DATA_VALID_DEL13__0,
    load_CRC8,
    start_CRC8,
    txstatplus_int0_out,
    append_end_frame,
    \TX_DATA_DEL14_reg[32]_0 ,
    \TX_DATA_DEL14_reg[18] ,
    \TX_DATA_DEL14_reg[18]_0 ,
    \TX_DATA_DEL14_reg[58]_0 ,
    \TX_DATA_DEL14_reg[58]_1 ,
    \TX_DATA_DEL14_reg[57] ,
    \TX_DATA_DEL14_reg[55] ,
    \TX_DATA_DEL14_reg[54] ,
    \TX_DATA_DEL14_reg[54]_0 ,
    \TX_DATA_DEL14_reg[53] ,
    \TX_DATA_DEL14_reg[52] ,
    \TX_DATA_DEL14_reg[51] ,
    \TX_DATA_DEL14_reg[49] ,
    \TX_DATA_DEL14_reg[49]_0 ,
    \TX_DATA_DEL14_reg[48] ,
    \TX_DATA_DEL14_reg[48]_0 ,
    \TX_DATA_DEL14_reg[39] ,
    \TX_DATA_DEL14_reg[38] ,
    \TX_DATA_DEL14_reg[33]_0 ,
    \TX_DATA_DEL14_reg[0] ,
    \TX_DATA_DEL14[57]_i_2_0 ,
    \TX_DATA_DEL14_reg[25] ,
    \TX_DATA_DEL14[57]_i_2_1 ,
    \TX_DATA_DEL14[63]_i_2_0 ,
    \TX_DATA_DEL14[57]_i_2_2 ,
    \TX_DATA_DEL14_reg[41] ,
    \TX_DATA_DEL14_reg[47] ,
    \CRC_OUT_reg[31]_0 ,
    \OVERFLOW_DATA_reg[19] ,
    clk_i,
    rst_i);
  output [23:0]D;
  output [0:0]E;
  output [63:0]\TX_DATA_VALID_DEL13_reg[7] ;
  input \TX_DATA_DEL14_reg[32] ;
  input fcs_enabled_int;
  input [0:0]TX_DATA_VALID_DEL13;
  input \TX_DATA_DEL14_reg[58] ;
  input [63:0]TX_DATA_DEL13;
  input \TX_DATA_DEL14_reg[50] ;
  input \TX_DATA_DEL14_reg[33] ;
  input \TX_DATA_DEL14_reg[26] ;
  input \OVERFLOW_DATA_reg[8] ;
  input \TX_DATA_DEL14_reg[21] ;
  input [7:0]Q;
  input \OVERFLOW_DATA_reg[2] ;
  input [0:0]txstatplus_int;
  input \OVERFLOW_DATA_reg[2]_0 ;
  input [5:0]TX_DATA_VALID_DEL13__0;
  input load_CRC8;
  input start_CRC8;
  input [0:0]txstatplus_int0_out;
  input append_end_frame;
  input \TX_DATA_DEL14_reg[32]_0 ;
  input \TX_DATA_DEL14_reg[18] ;
  input \TX_DATA_DEL14_reg[18]_0 ;
  input \TX_DATA_DEL14_reg[58]_0 ;
  input \TX_DATA_DEL14_reg[58]_1 ;
  input \TX_DATA_DEL14_reg[57] ;
  input \TX_DATA_DEL14_reg[55] ;
  input \TX_DATA_DEL14_reg[54] ;
  input \TX_DATA_DEL14_reg[54]_0 ;
  input \TX_DATA_DEL14_reg[53] ;
  input \TX_DATA_DEL14_reg[52] ;
  input \TX_DATA_DEL14_reg[51] ;
  input \TX_DATA_DEL14_reg[49] ;
  input \TX_DATA_DEL14_reg[49]_0 ;
  input \TX_DATA_DEL14_reg[48] ;
  input \TX_DATA_DEL14_reg[48]_0 ;
  input \TX_DATA_DEL14_reg[39] ;
  input [25:0]\TX_DATA_DEL14_reg[38] ;
  input \TX_DATA_DEL14_reg[33]_0 ;
  input \TX_DATA_DEL14_reg[0] ;
  input \TX_DATA_DEL14[57]_i_2_0 ;
  input \TX_DATA_DEL14_reg[25] ;
  input \TX_DATA_DEL14[57]_i_2_1 ;
  input \TX_DATA_DEL14[63]_i_2_0 ;
  input \TX_DATA_DEL14[57]_i_2_2 ;
  input \TX_DATA_DEL14_reg[41] ;
  input \TX_DATA_DEL14_reg[47] ;
  input [31:0]\CRC_OUT_reg[31]_0 ;
  input \OVERFLOW_DATA_reg[19] ;
  input clk_i;
  input rst_i;

  wire [31:0]CRC_OUT;
  wire \CRC_OUT[0]_i_1__2_n_0 ;
  wire \CRC_OUT[10]_i_1__2_n_0 ;
  wire \CRC_OUT[10]_i_2__2_n_0 ;
  wire \CRC_OUT[11]_i_1__2_n_0 ;
  wire \CRC_OUT[11]_i_2__2_n_0 ;
  wire \CRC_OUT[12]_i_1__2_n_0 ;
  wire \CRC_OUT[12]_i_2__2_n_0 ;
  wire \CRC_OUT[12]_i_3__1_n_0 ;
  wire \CRC_OUT[13]_i_1__2_n_0 ;
  wire \CRC_OUT[13]_i_2__2_n_0 ;
  wire \CRC_OUT[13]_i_3__2_n_0 ;
  wire \CRC_OUT[14]_i_1__2_n_0 ;
  wire \CRC_OUT[14]_i_2__1_n_0 ;
  wire \CRC_OUT[14]_i_3__2_n_0 ;
  wire \CRC_OUT[14]_i_4__1_n_0 ;
  wire \CRC_OUT[15]_i_1__2_n_0 ;
  wire \CRC_OUT[15]_i_2__2_n_0 ;
  wire \CRC_OUT[15]_i_3__2_n_0 ;
  wire \CRC_OUT[16]_i_1__2_n_0 ;
  wire \CRC_OUT[16]_i_2__2_n_0 ;
  wire \CRC_OUT[16]_i_3__2_n_0 ;
  wire \CRC_OUT[16]_i_4__2_n_0 ;
  wire \CRC_OUT[17]_i_1__2_n_0 ;
  wire \CRC_OUT[17]_i_2__2_n_0 ;
  wire \CRC_OUT[17]_i_3__1_n_0 ;
  wire \CRC_OUT[18]_i_1__2_n_0 ;
  wire \CRC_OUT[18]_i_2__2_n_0 ;
  wire \CRC_OUT[19]_i_1__2_n_0 ;
  wire \CRC_OUT[19]_i_2__2_n_0 ;
  wire \CRC_OUT[1]_i_1__2_n_0 ;
  wire \CRC_OUT[20]_i_1__2_n_0 ;
  wire \CRC_OUT[21]_i_1__2_n_0 ;
  wire \CRC_OUT[22]_i_1__2_n_0 ;
  wire \CRC_OUT[23]_i_1__2_n_0 ;
  wire \CRC_OUT[23]_i_2__2_n_0 ;
  wire \CRC_OUT[24]_i_1__2_n_0 ;
  wire \CRC_OUT[24]_i_2__2_n_0 ;
  wire \CRC_OUT[24]_i_3__2_n_0 ;
  wire \CRC_OUT[25]_i_1__2_n_0 ;
  wire \CRC_OUT[25]_i_2__2_n_0 ;
  wire \CRC_OUT[26]_i_1__2_n_0 ;
  wire \CRC_OUT[26]_i_2__2_n_0 ;
  wire \CRC_OUT[27]_i_1__2_n_0 ;
  wire \CRC_OUT[27]_i_2__2_n_0 ;
  wire \CRC_OUT[27]_i_3__1_n_0 ;
  wire \CRC_OUT[27]_i_4__1_n_0 ;
  wire \CRC_OUT[28]_i_1__2_n_0 ;
  wire \CRC_OUT[28]_i_2__2_n_0 ;
  wire \CRC_OUT[29]_i_1__2_n_0 ;
  wire \CRC_OUT[29]_i_2__2_n_0 ;
  wire \CRC_OUT[2]_i_1__2_n_0 ;
  wire \CRC_OUT[2]_i_2__2_n_0 ;
  wire \CRC_OUT[30]_i_1__2_n_0 ;
  wire \CRC_OUT[30]_i_2__2_n_0 ;
  wire \CRC_OUT[31]_i_2__1_n_0 ;
  wire \CRC_OUT[3]_i_1__2_n_0 ;
  wire \CRC_OUT[3]_i_2__1_n_0 ;
  wire \CRC_OUT[4]_i_1__2_n_0 ;
  wire \CRC_OUT[4]_i_2__2_n_0 ;
  wire \CRC_OUT[4]_i_3__1_n_0 ;
  wire \CRC_OUT[5]_i_1__2_n_0 ;
  wire \CRC_OUT[5]_i_2__2_n_0 ;
  wire \CRC_OUT[6]_i_1__2_n_0 ;
  wire \CRC_OUT[6]_i_2__2_n_0 ;
  wire \CRC_OUT[7]_i_1__2_n_0 ;
  wire \CRC_OUT[7]_i_2__2_n_0 ;
  wire \CRC_OUT[7]_i_3__1_n_0 ;
  wire \CRC_OUT[8]_i_1__2_n_0 ;
  wire \CRC_OUT[9]_i_1__2_n_0 ;
  wire \CRC_OUT[9]_i_2__2_n_0 ;
  wire [31:0]\CRC_OUT_reg[31]_0 ;
  wire [23:0]D;
  wire [0:0]E;
  wire \OVERFLOW_DATA[0]_i_2_n_0 ;
  wire \OVERFLOW_DATA[11]_i_2_n_0 ;
  wire \OVERFLOW_DATA[12]_i_2_n_0 ;
  wire \OVERFLOW_DATA[13]_i_2_n_0 ;
  wire \OVERFLOW_DATA[14]_i_2_n_0 ;
  wire \OVERFLOW_DATA[15]_i_2_n_0 ;
  wire \OVERFLOW_DATA[1]_i_2_n_0 ;
  wire \OVERFLOW_DATA[1]_i_3_n_0 ;
  wire \OVERFLOW_DATA[2]_i_2_n_0 ;
  wire \OVERFLOW_DATA[2]_i_3_n_0 ;
  wire \OVERFLOW_DATA[3]_i_2_n_0 ;
  wire \OVERFLOW_DATA[4]_i_2_n_0 ;
  wire \OVERFLOW_DATA[5]_i_2_n_0 ;
  wire \OVERFLOW_DATA[6]_i_2_n_0 ;
  wire \OVERFLOW_DATA[7]_i_2_n_0 ;
  wire \OVERFLOW_DATA[8]_i_3_n_0 ;
  wire \OVERFLOW_DATA[9]_i_2_n_0 ;
  wire \OVERFLOW_DATA_reg[19] ;
  wire \OVERFLOW_DATA_reg[2] ;
  wire \OVERFLOW_DATA_reg[2]_0 ;
  wire \OVERFLOW_DATA_reg[8] ;
  wire [7:0]Q;
  wire [63:0]TX_DATA_DEL13;
  wire \TX_DATA_DEL14[0]_i_2_n_0 ;
  wire \TX_DATA_DEL14[11]_i_2_n_0 ;
  wire \TX_DATA_DEL14[12]_i_2_n_0 ;
  wire \TX_DATA_DEL14[13]_i_2_n_0 ;
  wire \TX_DATA_DEL14[14]_i_2_n_0 ;
  wire \TX_DATA_DEL14[15]_i_3_n_0 ;
  wire \TX_DATA_DEL14[16]_i_2_n_0 ;
  wire \TX_DATA_DEL14[17]_i_2_n_0 ;
  wire \TX_DATA_DEL14[18]_i_2_n_0 ;
  wire \TX_DATA_DEL14[18]_i_3_n_0 ;
  wire \TX_DATA_DEL14[19]_i_2_n_0 ;
  wire \TX_DATA_DEL14[1]_i_2_n_0 ;
  wire \TX_DATA_DEL14[20]_i_2_n_0 ;
  wire \TX_DATA_DEL14[21]_i_2_n_0 ;
  wire \TX_DATA_DEL14[22]_i_2_n_0 ;
  wire \TX_DATA_DEL14[23]_i_3_n_0 ;
  wire \TX_DATA_DEL14[24]_i_2_n_0 ;
  wire \TX_DATA_DEL14[24]_i_3_n_0 ;
  wire \TX_DATA_DEL14[25]_i_2_n_0 ;
  wire \TX_DATA_DEL14[25]_i_3_n_0 ;
  wire \TX_DATA_DEL14[26]_i_2_n_0 ;
  wire \TX_DATA_DEL14[26]_i_3_n_0 ;
  wire \TX_DATA_DEL14[27]_i_2_n_0 ;
  wire \TX_DATA_DEL14[27]_i_3_n_0 ;
  wire \TX_DATA_DEL14[27]_i_4_n_0 ;
  wire \TX_DATA_DEL14[27]_i_5_n_0 ;
  wire \TX_DATA_DEL14[28]_i_2_n_0 ;
  wire \TX_DATA_DEL14[28]_i_3_n_0 ;
  wire \TX_DATA_DEL14[28]_i_4_n_0 ;
  wire \TX_DATA_DEL14[28]_i_5_n_0 ;
  wire \TX_DATA_DEL14[29]_i_2_n_0 ;
  wire \TX_DATA_DEL14[29]_i_3_n_0 ;
  wire \TX_DATA_DEL14[29]_i_4_n_0 ;
  wire \TX_DATA_DEL14[29]_i_5_n_0 ;
  wire \TX_DATA_DEL14[2]_i_2_n_0 ;
  wire \TX_DATA_DEL14[30]_i_2_n_0 ;
  wire \TX_DATA_DEL14[30]_i_3_n_0 ;
  wire \TX_DATA_DEL14[30]_i_4_n_0 ;
  wire \TX_DATA_DEL14[30]_i_5_n_0 ;
  wire \TX_DATA_DEL14[31]_i_2_n_0 ;
  wire \TX_DATA_DEL14[31]_i_3_n_0 ;
  wire \TX_DATA_DEL14[31]_i_4_n_0 ;
  wire \TX_DATA_DEL14[31]_i_5_n_0 ;
  wire \TX_DATA_DEL14[32]_i_2_n_0 ;
  wire \TX_DATA_DEL14[32]_i_3_n_0 ;
  wire \TX_DATA_DEL14[33]_i_2_n_0 ;
  wire \TX_DATA_DEL14[33]_i_3_n_0 ;
  wire \TX_DATA_DEL14[33]_i_5_n_0 ;
  wire \TX_DATA_DEL14[34]_i_2_n_0 ;
  wire \TX_DATA_DEL14[34]_i_3_n_0 ;
  wire \TX_DATA_DEL14[35]_i_2_n_0 ;
  wire \TX_DATA_DEL14[35]_i_3_n_0 ;
  wire \TX_DATA_DEL14[36]_i_2_n_0 ;
  wire \TX_DATA_DEL14[36]_i_3_n_0 ;
  wire \TX_DATA_DEL14[36]_i_4_n_0 ;
  wire \TX_DATA_DEL14[37]_i_2_n_0 ;
  wire \TX_DATA_DEL14[37]_i_3_n_0 ;
  wire \TX_DATA_DEL14[37]_i_4_n_0 ;
  wire \TX_DATA_DEL14[38]_i_2_n_0 ;
  wire \TX_DATA_DEL14[38]_i_3_n_0 ;
  wire \TX_DATA_DEL14[39]_i_2_n_0 ;
  wire \TX_DATA_DEL14[39]_i_4_n_0 ;
  wire \TX_DATA_DEL14[39]_i_6_n_0 ;
  wire \TX_DATA_DEL14[3]_i_2_n_0 ;
  wire \TX_DATA_DEL14[40]_i_2_n_0 ;
  wire \TX_DATA_DEL14[40]_i_3_n_0 ;
  wire \TX_DATA_DEL14[41]_i_2_n_0 ;
  wire \TX_DATA_DEL14[41]_i_3_n_0 ;
  wire \TX_DATA_DEL14[41]_i_4_n_0 ;
  wire \TX_DATA_DEL14[42]_i_2_n_0 ;
  wire \TX_DATA_DEL14[42]_i_3_n_0 ;
  wire \TX_DATA_DEL14[42]_i_4_n_0 ;
  wire \TX_DATA_DEL14[43]_i_2_n_0 ;
  wire \TX_DATA_DEL14[43]_i_3_n_0 ;
  wire \TX_DATA_DEL14[43]_i_4_n_0 ;
  wire \TX_DATA_DEL14[44]_i_2_n_0 ;
  wire \TX_DATA_DEL14[44]_i_3_n_0 ;
  wire \TX_DATA_DEL14[45]_i_2_n_0 ;
  wire \TX_DATA_DEL14[45]_i_3_n_0 ;
  wire \TX_DATA_DEL14[46]_i_2_n_0 ;
  wire \TX_DATA_DEL14[46]_i_3_n_0 ;
  wire \TX_DATA_DEL14[46]_i_4_n_0 ;
  wire \TX_DATA_DEL14[47]_i_2_n_0 ;
  wire \TX_DATA_DEL14[47]_i_4_n_0 ;
  wire \TX_DATA_DEL14[48]_i_2_n_0 ;
  wire \TX_DATA_DEL14[48]_i_3_n_0 ;
  wire \TX_DATA_DEL14[48]_i_4_n_0 ;
  wire \TX_DATA_DEL14[49]_i_2_n_0 ;
  wire \TX_DATA_DEL14[49]_i_3_n_0 ;
  wire \TX_DATA_DEL14[49]_i_4_n_0 ;
  wire \TX_DATA_DEL14[4]_i_2_n_0 ;
  wire \TX_DATA_DEL14[50]_i_2_n_0 ;
  wire \TX_DATA_DEL14[50]_i_4_n_0 ;
  wire \TX_DATA_DEL14[51]_i_2_n_0 ;
  wire \TX_DATA_DEL14[51]_i_3_n_0 ;
  wire \TX_DATA_DEL14[51]_i_4_n_0 ;
  wire \TX_DATA_DEL14[51]_i_6_n_0 ;
  wire \TX_DATA_DEL14[52]_i_2_n_0 ;
  wire \TX_DATA_DEL14[52]_i_4_n_0 ;
  wire \TX_DATA_DEL14[52]_i_5_n_0 ;
  wire \TX_DATA_DEL14[53]_i_2_n_0 ;
  wire \TX_DATA_DEL14[53]_i_4_n_0 ;
  wire \TX_DATA_DEL14[53]_i_5_n_0 ;
  wire \TX_DATA_DEL14[54]_i_2_n_0 ;
  wire \TX_DATA_DEL14[54]_i_3_n_0 ;
  wire \TX_DATA_DEL14[54]_i_4_n_0 ;
  wire \TX_DATA_DEL14[54]_i_7_n_0 ;
  wire \TX_DATA_DEL14[55]_i_2_n_0 ;
  wire \TX_DATA_DEL14[55]_i_4_n_0 ;
  wire \TX_DATA_DEL14[55]_i_5_n_0 ;
  wire \TX_DATA_DEL14[56]_i_2_n_0 ;
  wire \TX_DATA_DEL14[56]_i_3_n_0 ;
  wire \TX_DATA_DEL14[56]_i_4_n_0 ;
  wire \TX_DATA_DEL14[56]_i_5_n_0 ;
  wire \TX_DATA_DEL14[56]_i_6_n_0 ;
  wire \TX_DATA_DEL14[57]_i_2_0 ;
  wire \TX_DATA_DEL14[57]_i_2_1 ;
  wire \TX_DATA_DEL14[57]_i_2_2 ;
  wire \TX_DATA_DEL14[57]_i_2_n_0 ;
  wire \TX_DATA_DEL14[57]_i_3_n_0 ;
  wire \TX_DATA_DEL14[57]_i_4_n_0 ;
  wire \TX_DATA_DEL14[57]_i_5_n_0 ;
  wire \TX_DATA_DEL14[58]_i_2_n_0 ;
  wire \TX_DATA_DEL14[58]_i_4_n_0 ;
  wire \TX_DATA_DEL14[59]_i_2_n_0 ;
  wire \TX_DATA_DEL14[59]_i_3_n_0 ;
  wire \TX_DATA_DEL14[59]_i_4_n_0 ;
  wire \TX_DATA_DEL14[5]_i_2_n_0 ;
  wire \TX_DATA_DEL14[60]_i_2_n_0 ;
  wire \TX_DATA_DEL14[60]_i_3_n_0 ;
  wire \TX_DATA_DEL14[60]_i_4_n_0 ;
  wire \TX_DATA_DEL14[61]_i_2_n_0 ;
  wire \TX_DATA_DEL14[61]_i_3_n_0 ;
  wire \TX_DATA_DEL14[61]_i_4_n_0 ;
  wire \TX_DATA_DEL14[62]_i_2_n_0 ;
  wire \TX_DATA_DEL14[62]_i_3_n_0 ;
  wire \TX_DATA_DEL14[62]_i_4_n_0 ;
  wire \TX_DATA_DEL14[63]_i_2_0 ;
  wire \TX_DATA_DEL14[63]_i_2_n_0 ;
  wire \TX_DATA_DEL14[63]_i_3_n_0 ;
  wire \TX_DATA_DEL14[63]_i_6_n_0 ;
  wire \TX_DATA_DEL14[6]_i_2_n_0 ;
  wire \TX_DATA_DEL14[7]_i_2_n_0 ;
  wire \TX_DATA_DEL14[8]_i_2_n_0 ;
  wire \TX_DATA_DEL14[9]_i_2_n_0 ;
  wire \TX_DATA_DEL14_reg[0] ;
  wire \TX_DATA_DEL14_reg[18] ;
  wire \TX_DATA_DEL14_reg[18]_0 ;
  wire \TX_DATA_DEL14_reg[21] ;
  wire \TX_DATA_DEL14_reg[25] ;
  wire \TX_DATA_DEL14_reg[26] ;
  wire \TX_DATA_DEL14_reg[32] ;
  wire \TX_DATA_DEL14_reg[32]_0 ;
  wire \TX_DATA_DEL14_reg[33] ;
  wire \TX_DATA_DEL14_reg[33]_0 ;
  wire [25:0]\TX_DATA_DEL14_reg[38] ;
  wire \TX_DATA_DEL14_reg[39] ;
  wire \TX_DATA_DEL14_reg[41] ;
  wire \TX_DATA_DEL14_reg[47] ;
  wire \TX_DATA_DEL14_reg[48] ;
  wire \TX_DATA_DEL14_reg[48]_0 ;
  wire \TX_DATA_DEL14_reg[49] ;
  wire \TX_DATA_DEL14_reg[49]_0 ;
  wire \TX_DATA_DEL14_reg[50] ;
  wire \TX_DATA_DEL14_reg[51] ;
  wire \TX_DATA_DEL14_reg[52] ;
  wire \TX_DATA_DEL14_reg[53] ;
  wire \TX_DATA_DEL14_reg[54] ;
  wire \TX_DATA_DEL14_reg[54]_0 ;
  wire \TX_DATA_DEL14_reg[55] ;
  wire \TX_DATA_DEL14_reg[57] ;
  wire \TX_DATA_DEL14_reg[58] ;
  wire \TX_DATA_DEL14_reg[58]_0 ;
  wire \TX_DATA_DEL14_reg[58]_1 ;
  wire [0:0]TX_DATA_VALID_DEL13;
  wire [5:0]TX_DATA_VALID_DEL13__0;
  wire [63:0]\TX_DATA_VALID_DEL13_reg[7] ;
  wire append_end_frame;
  wire clk_i;
  wire fcs_enabled_int;
  wire load_CRC8;
  wire rst_i;
  wire start_CRC8;
  wire [0:0]txstatplus_int;
  wire [0:0]txstatplus_int0_out;

  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[0]_i_1__2 
       (.I0(CRC_OUT[24]),
        .I1(Q[0]),
        .I2(Q[6]),
        .I3(CRC_OUT[30]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [0]),
        .O(\CRC_OUT[0]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[10]_i_1__2 
       (.I0(CRC_OUT[26]),
        .I1(CRC_OUT[2]),
        .I2(\CRC_OUT[14]_i_4__1_n_0 ),
        .I3(\CRC_OUT[10]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [10]),
        .O(\CRC_OUT[10]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair385" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \CRC_OUT[10]_i_2__2 
       (.I0(Q[5]),
        .I1(CRC_OUT[29]),
        .I2(Q[0]),
        .I3(CRC_OUT[24]),
        .I4(Q[2]),
        .O(\CRC_OUT[10]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair391" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \CRC_OUT[11]_i_1__2 
       (.I0(CRC_OUT[3]),
        .I1(\CRC_OUT[11]_i_2__2_n_0 ),
        .I2(start_CRC8),
        .I3(\CRC_OUT_reg[31]_0 [11]),
        .O(\CRC_OUT[11]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair376" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[11]_i_2__2 
       (.I0(CRC_OUT[27]),
        .I1(Q[3]),
        .I2(CRC_OUT[28]),
        .I3(Q[4]),
        .I4(\CRC_OUT[12]_i_2__2_n_0 ),
        .O(\CRC_OUT[11]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[12]_i_1__2 
       (.I0(\CRC_OUT[12]_i_2__2_n_0 ),
        .I1(CRC_OUT[30]),
        .I2(\CRC_OUT[24]_i_3__2_n_0 ),
        .I3(\CRC_OUT[12]_i_3__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [12]),
        .O(\CRC_OUT[12]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair387" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[12]_i_2__2 
       (.I0(Q[1]),
        .I1(CRC_OUT[25]),
        .I2(CRC_OUT[24]),
        .I3(Q[0]),
        .O(\CRC_OUT[12]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[12]_i_3__1 
       (.I0(CRC_OUT[28]),
        .I1(CRC_OUT[29]),
        .I2(Q[4]),
        .I3(CRC_OUT[4]),
        .I4(Q[5]),
        .I5(Q[6]),
        .O(\CRC_OUT[12]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[13]_i_1__2 
       (.I0(\CRC_OUT[13]_i_2__2_n_0 ),
        .I1(CRC_OUT[27]),
        .I2(CRC_OUT[26]),
        .I3(\CRC_OUT[13]_i_3__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [13]),
        .O(\CRC_OUT[13]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair393" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \CRC_OUT[13]_i_2__2 
       (.I0(CRC_OUT[30]),
        .I1(CRC_OUT[31]),
        .I2(CRC_OUT[29]),
        .O(\CRC_OUT[13]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_3__2 
       (.I0(Q[2]),
        .I1(CRC_OUT[5]),
        .I2(\CRC_OUT[27]_i_2__2_n_0 ),
        .I3(\CRC_OUT[19]_i_2__2_n_0 ),
        .I4(Q[5]),
        .I5(Q[6]),
        .O(\CRC_OUT[13]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[14]_i_1__2 
       (.I0(\CRC_OUT[14]_i_2__1_n_0 ),
        .I1(CRC_OUT[6]),
        .I2(\CRC_OUT[14]_i_3__2_n_0 ),
        .I3(\CRC_OUT[14]_i_4__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [14]),
        .O(\CRC_OUT[14]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[14]_i_2__1 
       (.I0(Q[2]),
        .I1(CRC_OUT[26]),
        .I2(CRC_OUT[30]),
        .I3(CRC_OUT[28]),
        .I4(Q[4]),
        .I5(CRC_OUT[31]),
        .O(\CRC_OUT[14]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair389" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[14]_i_3__2 
       (.I0(Q[7]),
        .I1(Q[6]),
        .O(\CRC_OUT[14]_i_3__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair376" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \CRC_OUT[14]_i_4__1 
       (.I0(CRC_OUT[27]),
        .I1(Q[3]),
        .O(\CRC_OUT[14]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[15]_i_1__2 
       (.I0(\CRC_OUT[15]_i_2__2_n_0 ),
        .I1(\CRC_OUT[15]_i_3__2_n_0 ),
        .I2(CRC_OUT[29]),
        .I3(CRC_OUT[31]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [15]),
        .O(\CRC_OUT[15]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair372" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[15]_i_2__2 
       (.I0(Q[7]),
        .I1(Q[5]),
        .I2(Q[4]),
        .I3(CRC_OUT[7]),
        .I4(Q[3]),
        .O(\CRC_OUT[15]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair400" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[15]_i_3__2 
       (.I0(CRC_OUT[28]),
        .I1(CRC_OUT[27]),
        .O(\CRC_OUT[15]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[16]_i_1__2 
       (.I0(\CRC_OUT[16]_i_2__2_n_0 ),
        .I1(\CRC_OUT[16]_i_3__2_n_0 ),
        .I2(\CRC_OUT[16]_i_4__2_n_0 ),
        .I3(CRC_OUT[8]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [16]),
        .O(\CRC_OUT[16]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair380" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[16]_i_2__2 
       (.I0(Q[0]),
        .I1(CRC_OUT[24]),
        .O(\CRC_OUT[16]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair399" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \CRC_OUT[16]_i_3__2 
       (.I0(CRC_OUT[29]),
        .I1(CRC_OUT[28]),
        .O(\CRC_OUT[16]_i_3__2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \CRC_OUT[16]_i_4__2 
       (.I0(Q[5]),
        .I1(Q[4]),
        .O(\CRC_OUT[16]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[17]_i_1__2 
       (.I0(\CRC_OUT[17]_i_2__2_n_0 ),
        .I1(Q[6]),
        .I2(CRC_OUT[9]),
        .I3(\CRC_OUT[17]_i_3__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [17]),
        .O(\CRC_OUT[17]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair387" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \CRC_OUT[17]_i_2__2 
       (.I0(CRC_OUT[30]),
        .I1(Q[1]),
        .I2(CRC_OUT[25]),
        .O(\CRC_OUT[17]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair379" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_3__1 
       (.I0(CRC_OUT[29]),
        .I1(Q[5]),
        .O(\CRC_OUT[17]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[18]_i_1__2 
       (.I0(CRC_OUT[31]),
        .I1(CRC_OUT[26]),
        .I2(CRC_OUT[10]),
        .I3(\CRC_OUT[18]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [18]),
        .O(\CRC_OUT[18]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair392" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[18]_i_2__2 
       (.I0(Q[6]),
        .I1(Q[7]),
        .I2(Q[2]),
        .I3(CRC_OUT[30]),
        .O(\CRC_OUT[18]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[19]_i_1__2 
       (.I0(CRC_OUT[27]),
        .I1(CRC_OUT[31]),
        .I2(\CRC_OUT[19]_i_2__2_n_0 ),
        .I3(CRC_OUT[11]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [19]),
        .O(\CRC_OUT[19]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair404" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[19]_i_2__2 
       (.I0(Q[7]),
        .I1(Q[3]),
        .O(\CRC_OUT[19]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[1]_i_1__2 
       (.I0(\CRC_OUT[12]_i_2__2_n_0 ),
        .I1(CRC_OUT[30]),
        .I2(Q[6]),
        .I3(\CRC_OUT[24]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [1]),
        .O(\CRC_OUT[1]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair384" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[20]_i_1__2 
       (.I0(CRC_OUT[12]),
        .I1(Q[4]),
        .I2(CRC_OUT[28]),
        .I3(start_CRC8),
        .I4(\CRC_OUT_reg[31]_0 [20]),
        .O(\CRC_OUT[20]_i_1__2_n_0 ));
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[21]_i_1__2 
       (.I0(CRC_OUT[13]),
        .I1(Q[5]),
        .I2(CRC_OUT[29]),
        .I3(start_CRC8),
        .I4(\CRC_OUT_reg[31]_0 [21]),
        .O(\CRC_OUT[21]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair380" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[22]_i_1__2 
       (.I0(CRC_OUT[14]),
        .I1(CRC_OUT[24]),
        .I2(Q[0]),
        .I3(start_CRC8),
        .I4(\CRC_OUT_reg[31]_0 [22]),
        .O(\CRC_OUT[22]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[23]_i_1__2 
       (.I0(CRC_OUT[25]),
        .I1(Q[1]),
        .I2(CRC_OUT[15]),
        .I3(\CRC_OUT[23]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [23]),
        .O(\CRC_OUT[23]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair386" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[23]_i_2__2 
       (.I0(CRC_OUT[24]),
        .I1(Q[0]),
        .I2(Q[6]),
        .I3(CRC_OUT[30]),
        .O(\CRC_OUT[23]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[24]_i_1__2 
       (.I0(\CRC_OUT[24]_i_2__2_n_0 ),
        .I1(CRC_OUT[16]),
        .I2(\CRC_OUT[24]_i_3__2_n_0 ),
        .I3(\CRC_OUT[27]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [24]),
        .O(\CRC_OUT[24]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair392" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_2__2 
       (.I0(CRC_OUT[31]),
        .I1(Q[7]),
        .O(\CRC_OUT[24]_i_2__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_3__2 
       (.I0(Q[2]),
        .I1(CRC_OUT[26]),
        .O(\CRC_OUT[24]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[25]_i_1__2 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(\CRC_OUT[25]_i_2__2_n_0 ),
        .I3(CRC_OUT[17]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [25]),
        .O(\CRC_OUT[25]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair400" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \CRC_OUT[25]_i_2__2 
       (.I0(CRC_OUT[27]),
        .I1(CRC_OUT[26]),
        .O(\CRC_OUT[25]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[26]_i_1__2 
       (.I0(Q[0]),
        .I1(CRC_OUT[24]),
        .I2(CRC_OUT[30]),
        .I3(\CRC_OUT[26]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [26]),
        .O(\CRC_OUT[26]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[26]_i_2__2 
       (.I0(Q[4]),
        .I1(Q[3]),
        .I2(Q[6]),
        .I3(CRC_OUT[28]),
        .I4(CRC_OUT[27]),
        .I5(CRC_OUT[18]),
        .O(\CRC_OUT[26]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[27]_i_1__2 
       (.I0(\CRC_OUT[27]_i_2__2_n_0 ),
        .I1(\CRC_OUT[27]_i_3__1_n_0 ),
        .I2(\CRC_OUT[27]_i_4__1_n_0 ),
        .I3(CRC_OUT[19]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [27]),
        .O(\CRC_OUT[27]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair388" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[27]_i_2__2 
       (.I0(CRC_OUT[25]),
        .I1(Q[1]),
        .O(\CRC_OUT[27]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair393" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[27]_i_3__1 
       (.I0(CRC_OUT[28]),
        .I1(CRC_OUT[31]),
        .I2(CRC_OUT[29]),
        .O(\CRC_OUT[27]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair372" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[27]_i_4__1 
       (.I0(Q[4]),
        .I1(Q[5]),
        .I2(Q[7]),
        .O(\CRC_OUT[27]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[28]_i_1__2 
       (.I0(CRC_OUT[29]),
        .I1(Q[2]),
        .I2(CRC_OUT[20]),
        .I3(\CRC_OUT[28]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [28]),
        .O(\CRC_OUT[28]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair389" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_2__2 
       (.I0(Q[6]),
        .I1(Q[5]),
        .I2(CRC_OUT[26]),
        .I3(CRC_OUT[30]),
        .O(\CRC_OUT[28]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[29]_i_1__2 
       (.I0(Q[7]),
        .I1(Q[6]),
        .I2(CRC_OUT[21]),
        .I3(\CRC_OUT[29]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [29]),
        .O(\CRC_OUT[29]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair390" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[29]_i_2__2 
       (.I0(CRC_OUT[27]),
        .I1(CRC_OUT[31]),
        .I2(Q[3]),
        .I3(CRC_OUT[30]),
        .O(\CRC_OUT[29]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[2]_i_1__2 
       (.I0(CRC_OUT[31]),
        .I1(CRC_OUT[26]),
        .I2(\CRC_OUT[14]_i_3__2_n_0 ),
        .I3(\CRC_OUT[2]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [2]),
        .O(\CRC_OUT[2]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[2]_i_2__2 
       (.I0(CRC_OUT[25]),
        .I1(Q[1]),
        .I2(CRC_OUT[30]),
        .I3(Q[0]),
        .I4(CRC_OUT[24]),
        .I5(Q[2]),
        .O(\CRC_OUT[2]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[30]_i_1__2 
       (.I0(Q[7]),
        .I1(CRC_OUT[31]),
        .I2(\CRC_OUT[30]_i_2__2_n_0 ),
        .I3(CRC_OUT[22]),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [30]),
        .O(\CRC_OUT[30]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair384" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[30]_i_2__2 
       (.I0(CRC_OUT[28]),
        .I1(Q[4]),
        .O(\CRC_OUT[30]_i_2__2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \CRC_OUT[31]_i_1__0 
       (.I0(load_CRC8),
        .I1(start_CRC8),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair379" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[31]_i_2__1 
       (.I0(CRC_OUT[23]),
        .I1(Q[5]),
        .I2(CRC_OUT[29]),
        .I3(start_CRC8),
        .I4(\CRC_OUT_reg[31]_0 [31]),
        .O(\CRC_OUT[31]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[3]_i_1__2 
       (.I0(\CRC_OUT[19]_i_2__2_n_0 ),
        .I1(\CRC_OUT[27]_i_2__2_n_0 ),
        .I2(\CRC_OUT[24]_i_3__2_n_0 ),
        .I3(\CRC_OUT[3]_i_2__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [3]),
        .O(\CRC_OUT[3]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair390" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[3]_i_2__1 
       (.I0(CRC_OUT[31]),
        .I1(CRC_OUT[27]),
        .O(\CRC_OUT[3]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[4]_i_1__2 
       (.I0(\CRC_OUT[4]_i_2__2_n_0 ),
        .I1(CRC_OUT[28]),
        .I2(CRC_OUT[27]),
        .I3(\CRC_OUT[4]_i_3__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [4]),
        .O(\CRC_OUT[4]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair385" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[4]_i_2__2 
       (.I0(Q[2]),
        .I1(CRC_OUT[24]),
        .I2(Q[0]),
        .O(\CRC_OUT[4]_i_2__2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[4]_i_3__1 
       (.I0(CRC_OUT[26]),
        .I1(CRC_OUT[30]),
        .I2(Q[4]),
        .I3(Q[3]),
        .I4(Q[6]),
        .O(\CRC_OUT[4]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[5]_i_1__2 
       (.I0(\CRC_OUT[13]_i_2__2_n_0 ),
        .I1(CRC_OUT[28]),
        .I2(CRC_OUT[27]),
        .I3(\CRC_OUT[5]_i_2__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [5]),
        .O(\CRC_OUT[5]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[5]_i_2__2 
       (.I0(\CRC_OUT[12]_i_2__2_n_0 ),
        .I1(Q[3]),
        .I2(Q[6]),
        .I3(Q[7]),
        .I4(Q[5]),
        .I5(Q[4]),
        .O(\CRC_OUT[5]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[6]_i_1__2 
       (.I0(\CRC_OUT[6]_i_2__2_n_0 ),
        .I1(CRC_OUT[30]),
        .I2(Q[2]),
        .I3(\CRC_OUT[27]_i_3__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [6]),
        .O(\CRC_OUT[6]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[6]_i_2__2 
       (.I0(Q[7]),
        .I1(Q[6]),
        .I2(CRC_OUT[26]),
        .I3(Q[5]),
        .I4(Q[4]),
        .I5(\CRC_OUT[27]_i_2__2_n_0 ),
        .O(\CRC_OUT[6]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[7]_i_1__2 
       (.I0(\CRC_OUT[7]_i_2__2_n_0 ),
        .I1(Q[5]),
        .I2(Q[7]),
        .I3(\CRC_OUT[7]_i_3__1_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [7]),
        .O(\CRC_OUT[7]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair404" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[7]_i_2__2 
       (.I0(Q[3]),
        .I1(Q[2]),
        .O(\CRC_OUT[7]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[7]_i_3__1 
       (.I0(CRC_OUT[26]),
        .I1(CRC_OUT[27]),
        .I2(Q[0]),
        .I3(CRC_OUT[24]),
        .I4(CRC_OUT[29]),
        .I5(CRC_OUT[31]),
        .O(\CRC_OUT[7]_i_3__1_n_0 ));
  LUT4 #(
    .INIT(16'h6F60)) 
    \CRC_OUT[8]_i_1__2 
       (.I0(CRC_OUT[0]),
        .I1(\CRC_OUT[11]_i_2__2_n_0 ),
        .I2(start_CRC8),
        .I3(\CRC_OUT_reg[31]_0 [8]),
        .O(\CRC_OUT[8]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[9]_i_1__2 
       (.I0(\CRC_OUT[9]_i_2__2_n_0 ),
        .I1(CRC_OUT[1]),
        .I2(\CRC_OUT[16]_i_3__2_n_0 ),
        .I3(\CRC_OUT[24]_i_3__2_n_0 ),
        .I4(start_CRC8),
        .I5(\CRC_OUT_reg[31]_0 [9]),
        .O(\CRC_OUT[9]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair388" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \CRC_OUT[9]_i_2__2 
       (.I0(Q[1]),
        .I1(CRC_OUT[25]),
        .I2(Q[4]),
        .I3(Q[5]),
        .O(\CRC_OUT[9]_i_2__2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[0]_i_1__2_n_0 ),
        .Q(CRC_OUT[0]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[10] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[10]_i_1__2_n_0 ),
        .Q(CRC_OUT[10]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[11] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[11]_i_1__2_n_0 ),
        .Q(CRC_OUT[11]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[12] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[12]_i_1__2_n_0 ),
        .Q(CRC_OUT[12]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[13] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[13]_i_1__2_n_0 ),
        .Q(CRC_OUT[13]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[14] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[14]_i_1__2_n_0 ),
        .Q(CRC_OUT[14]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[15] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[15]_i_1__2_n_0 ),
        .Q(CRC_OUT[15]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[16] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[16]_i_1__2_n_0 ),
        .Q(CRC_OUT[16]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[17] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[17]_i_1__2_n_0 ),
        .Q(CRC_OUT[17]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[18] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[18]_i_1__2_n_0 ),
        .Q(CRC_OUT[18]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[19] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[19]_i_1__2_n_0 ),
        .Q(CRC_OUT[19]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[1]_i_1__2_n_0 ),
        .Q(CRC_OUT[1]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[20] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[20]_i_1__2_n_0 ),
        .Q(CRC_OUT[20]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[21] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[21]_i_1__2_n_0 ),
        .Q(CRC_OUT[21]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[22] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[22]_i_1__2_n_0 ),
        .Q(CRC_OUT[22]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[23] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[23]_i_1__2_n_0 ),
        .Q(CRC_OUT[23]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[24] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[24]_i_1__2_n_0 ),
        .Q(CRC_OUT[24]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[25] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[25]_i_1__2_n_0 ),
        .Q(CRC_OUT[25]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[26] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[26]_i_1__2_n_0 ),
        .Q(CRC_OUT[26]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[27] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[27]_i_1__2_n_0 ),
        .Q(CRC_OUT[27]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[28] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[28]_i_1__2_n_0 ),
        .Q(CRC_OUT[28]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[29] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[29]_i_1__2_n_0 ),
        .Q(CRC_OUT[29]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[2]_i_1__2_n_0 ),
        .Q(CRC_OUT[2]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[30] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[30]_i_1__2_n_0 ),
        .Q(CRC_OUT[30]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[31] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[31]_i_2__1_n_0 ),
        .Q(CRC_OUT[31]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[3] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[3]_i_1__2_n_0 ),
        .Q(CRC_OUT[3]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[4] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[4]_i_1__2_n_0 ),
        .Q(CRC_OUT[4]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[5] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[5]_i_1__2_n_0 ),
        .Q(CRC_OUT[5]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[6] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[6]_i_1__2_n_0 ),
        .Q(CRC_OUT[6]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[7] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[7]_i_1__2_n_0 ),
        .Q(CRC_OUT[7]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[8] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[8]_i_1__2_n_0 ),
        .Q(CRC_OUT[8]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[9] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\CRC_OUT[9]_i_1__2_n_0 ),
        .Q(CRC_OUT[9]));
  LUT6 #(
    .INIT(64'h0000FFFFFF7FFF7F)) 
    \OVERFLOW_DATA[0]_i_1 
       (.I0(fcs_enabled_int),
        .I1(txstatplus_int),
        .I2(\OVERFLOW_DATA_reg[2]_0 ),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(\OVERFLOW_DATA[0]_i_2_n_0 ),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'h4070404040707373)) 
    \OVERFLOW_DATA[0]_i_2 
       (.I0(CRC_OUT[8]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[24]),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[16]),
        .O(\OVERFLOW_DATA[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFE0EFEFFFFFFFF)) 
    \OVERFLOW_DATA[10]_i_1 
       (.I0(\OVERFLOW_DATA_reg[2] ),
        .I1(CRC_OUT[26]),
        .I2(\OVERFLOW_DATA_reg[2]_0 ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[18]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[10]));
  LUT6 #(
    .INIT(64'h88888888B8888888)) 
    \OVERFLOW_DATA[11]_i_1 
       (.I0(\OVERFLOW_DATA[11]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[3]),
        .I2(fcs_enabled_int),
        .I3(txstatplus_int),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\OVERFLOW_DATA_reg[2] ),
        .O(D[11]));
  (* SOFT_HLUTNM = "soft_lutpair378" *) 
  LUT5 #(
    .INIT(32'hB0B3B080)) 
    \OVERFLOW_DATA[11]_i_2 
       (.I0(CRC_OUT[19]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(CRC_OUT[27]),
        .O(\OVERFLOW_DATA[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h88888888B8888888)) 
    \OVERFLOW_DATA[12]_i_1 
       (.I0(\OVERFLOW_DATA[12]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[3]),
        .I2(fcs_enabled_int),
        .I3(txstatplus_int),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\OVERFLOW_DATA_reg[2] ),
        .O(D[12]));
  (* SOFT_HLUTNM = "soft_lutpair381" *) 
  LUT5 #(
    .INIT(32'hB0B3B080)) 
    \OVERFLOW_DATA[12]_i_2 
       (.I0(CRC_OUT[20]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(CRC_OUT[28]),
        .O(\OVERFLOW_DATA[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h88888888B8888888)) 
    \OVERFLOW_DATA[13]_i_1 
       (.I0(\OVERFLOW_DATA[13]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[3]),
        .I2(fcs_enabled_int),
        .I3(txstatplus_int),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\OVERFLOW_DATA_reg[2] ),
        .O(D[13]));
  (* SOFT_HLUTNM = "soft_lutpair374" *) 
  LUT5 #(
    .INIT(32'hB0B3B080)) 
    \OVERFLOW_DATA[13]_i_2 
       (.I0(CRC_OUT[21]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(CRC_OUT[29]),
        .O(\OVERFLOW_DATA[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h88888888B8888888)) 
    \OVERFLOW_DATA[14]_i_1 
       (.I0(\OVERFLOW_DATA[14]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[3]),
        .I2(fcs_enabled_int),
        .I3(txstatplus_int),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\OVERFLOW_DATA_reg[2] ),
        .O(D[14]));
  (* SOFT_HLUTNM = "soft_lutpair375" *) 
  LUT5 #(
    .INIT(32'hB0B3B080)) 
    \OVERFLOW_DATA[14]_i_2 
       (.I0(CRC_OUT[22]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(CRC_OUT[30]),
        .O(\OVERFLOW_DATA[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h88888888B8888888)) 
    \OVERFLOW_DATA[15]_i_1 
       (.I0(\OVERFLOW_DATA[15]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[3]),
        .I2(fcs_enabled_int),
        .I3(txstatplus_int),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\OVERFLOW_DATA_reg[2] ),
        .O(D[15]));
  (* SOFT_HLUTNM = "soft_lutpair377" *) 
  LUT5 #(
    .INIT(32'hB0B3B080)) 
    \OVERFLOW_DATA[15]_i_2 
       (.I0(CRC_OUT[23]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(CRC_OUT[31]),
        .O(\OVERFLOW_DATA[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF55FFDFDFDFDF)) 
    \OVERFLOW_DATA[16]_i_1 
       (.I0(TX_DATA_VALID_DEL13__0[3]),
        .I1(\OVERFLOW_DATA_reg[2] ),
        .I2(txstatplus_int),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[24]),
        .I5(\OVERFLOW_DATA_reg[2]_0 ),
        .O(D[16]));
  LUT6 #(
    .INIT(64'hFF6E0F6EFFFFFFFF)) 
    \OVERFLOW_DATA[17]_i_1 
       (.I0(\OVERFLOW_DATA_reg[2] ),
        .I1(txstatplus_int),
        .I2(fcs_enabled_int),
        .I3(\OVERFLOW_DATA_reg[2]_0 ),
        .I4(CRC_OUT[25]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[17]));
  (* SOFT_HLUTNM = "soft_lutpair382" *) 
  LUT5 #(
    .INIT(32'hFF7FFFFF)) 
    \OVERFLOW_DATA[18]_i_1 
       (.I0(TX_DATA_VALID_DEL13__0[3]),
        .I1(TX_DATA_VALID_DEL13__0[5]),
        .I2(TX_DATA_VALID_DEL13__0[2]),
        .I3(CRC_OUT[26]),
        .I4(fcs_enabled_int),
        .O(D[18]));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \OVERFLOW_DATA[19]_i_1 
       (.I0(\OVERFLOW_DATA_reg[19] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[27]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[19]));
  LUT6 #(
    .INIT(64'h00000000FF6FFFFF)) 
    \OVERFLOW_DATA[1]_i_1 
       (.I0(\OVERFLOW_DATA_reg[2] ),
        .I1(txstatplus_int),
        .I2(TX_DATA_VALID_DEL13__0[2]),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(fcs_enabled_int),
        .I5(\OVERFLOW_DATA[1]_i_2_n_0 ),
        .O(D[1]));
  LUT6 #(
    .INIT(64'h00008B00FF008B00)) 
    \OVERFLOW_DATA[1]_i_2 
       (.I0(\OVERFLOW_DATA[1]_i_3_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2] ),
        .I2(CRC_OUT[17]),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\TX_DATA_DEL14[9]_i_2_n_0 ),
        .O(\OVERFLOW_DATA[1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair402" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \OVERFLOW_DATA[1]_i_3 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[25]),
        .O(\OVERFLOW_DATA[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \OVERFLOW_DATA[20]_i_1 
       (.I0(\OVERFLOW_DATA_reg[19] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[28]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[20]));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \OVERFLOW_DATA[21]_i_1 
       (.I0(\OVERFLOW_DATA_reg[19] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[29]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[21]));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \OVERFLOW_DATA[22]_i_1 
       (.I0(\OVERFLOW_DATA_reg[19] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[30]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[22]));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \OVERFLOW_DATA[23]_i_1 
       (.I0(\OVERFLOW_DATA_reg[19] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[31]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[23]));
  LUT6 #(
    .INIT(64'h00FF74FFFFFF74FF)) 
    \OVERFLOW_DATA[2]_i_1 
       (.I0(\OVERFLOW_DATA[2]_i_2_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2] ),
        .I2(CRC_OUT[18]),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(\OVERFLOW_DATA_reg[2]_0 ),
        .I5(\OVERFLOW_DATA[2]_i_3_n_0 ),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair382" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \OVERFLOW_DATA[2]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[26]),
        .O(\OVERFLOW_DATA[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair405" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \OVERFLOW_DATA[2]_i_3 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[10]),
        .O(\OVERFLOW_DATA[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808800008088)) 
    \OVERFLOW_DATA[3]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(txstatplus_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(TX_DATA_VALID_DEL13__0[3]),
        .I5(\OVERFLOW_DATA[3]_i_2_n_0 ),
        .O(D[3]));
  LUT6 #(
    .INIT(64'hB888BBBBB8888888)) 
    \OVERFLOW_DATA[3]_i_2 
       (.I0(\TX_DATA_DEL14[11]_i_2_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[27]),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[19]),
        .O(\OVERFLOW_DATA[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808800008088)) 
    \OVERFLOW_DATA[4]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(txstatplus_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(TX_DATA_VALID_DEL13__0[3]),
        .I5(\OVERFLOW_DATA[4]_i_2_n_0 ),
        .O(D[4]));
  LUT6 #(
    .INIT(64'hB888BBBBB8888888)) 
    \OVERFLOW_DATA[4]_i_2 
       (.I0(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[28]),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[20]),
        .O(\OVERFLOW_DATA[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808800008088)) 
    \OVERFLOW_DATA[5]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(txstatplus_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(TX_DATA_VALID_DEL13__0[3]),
        .I5(\OVERFLOW_DATA[5]_i_2_n_0 ),
        .O(D[5]));
  LUT6 #(
    .INIT(64'hB888BBBBB8888888)) 
    \OVERFLOW_DATA[5]_i_2 
       (.I0(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[29]),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[21]),
        .O(\OVERFLOW_DATA[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808800008088)) 
    \OVERFLOW_DATA[6]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(txstatplus_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(TX_DATA_VALID_DEL13__0[3]),
        .I5(\OVERFLOW_DATA[6]_i_2_n_0 ),
        .O(D[6]));
  LUT6 #(
    .INIT(64'hB888BBBBB8888888)) 
    \OVERFLOW_DATA[6]_i_2 
       (.I0(\TX_DATA_DEL14[14]_i_2_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[30]),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[22]),
        .O(\OVERFLOW_DATA[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808800008088)) 
    \OVERFLOW_DATA[7]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(txstatplus_int),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(TX_DATA_VALID_DEL13__0[3]),
        .I5(\OVERFLOW_DATA[7]_i_2_n_0 ),
        .O(D[7]));
  LUT6 #(
    .INIT(64'hB888BBBBB8888888)) 
    \OVERFLOW_DATA[7]_i_2 
       (.I0(\TX_DATA_DEL14[15]_i_3_n_0 ),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[31]),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[23]),
        .O(\OVERFLOW_DATA[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h002EFF2EFFFFFFFF)) 
    \OVERFLOW_DATA[8]_i_1 
       (.I0(CRC_OUT[24]),
        .I1(\OVERFLOW_DATA_reg[2] ),
        .I2(\OVERFLOW_DATA_reg[8] ),
        .I3(\OVERFLOW_DATA_reg[2]_0 ),
        .I4(\OVERFLOW_DATA[8]_i_3_n_0 ),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[8]));
  (* SOFT_HLUTNM = "soft_lutpair403" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \OVERFLOW_DATA[8]_i_3 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[16]),
        .O(\OVERFLOW_DATA[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFFF7FFF7F)) 
    \OVERFLOW_DATA[9]_i_1 
       (.I0(fcs_enabled_int),
        .I1(txstatplus_int),
        .I2(\OVERFLOW_DATA_reg[2]_0 ),
        .I3(\OVERFLOW_DATA_reg[2] ),
        .I4(\OVERFLOW_DATA[9]_i_2_n_0 ),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(D[9]));
  LUT6 #(
    .INIT(64'h4070404040707373)) 
    \OVERFLOW_DATA[9]_i_2 
       (.I0(CRC_OUT[17]),
        .I1(\OVERFLOW_DATA_reg[2]_0 ),
        .I2(fcs_enabled_int),
        .I3(txstatplus_int),
        .I4(\OVERFLOW_DATA_reg[2] ),
        .I5(CRC_OUT[25]),
        .O(\OVERFLOW_DATA[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[0]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [0]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[0]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [0]));
  (* SOFT_HLUTNM = "soft_lutpair398" *) 
  LUT3 #(
    .INIT(8'hC5)) 
    \TX_DATA_DEL14[0]_i_2 
       (.I0(txstatplus_int),
        .I1(CRC_OUT[0]),
        .I2(fcs_enabled_int),
        .O(\TX_DATA_DEL14[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB00F08888)) 
    \TX_DATA_DEL14[10]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [10]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(\OVERFLOW_DATA[2]_i_3_n_0 ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[10]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [10]));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[11]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [11]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[11]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[11]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [11]));
  (* SOFT_HLUTNM = "soft_lutpair398" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[11]_i_2 
       (.I0(CRC_OUT[11]),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .O(\TX_DATA_DEL14[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[12]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [12]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[12]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [12]));
  (* SOFT_HLUTNM = "soft_lutpair397" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[12]_i_2 
       (.I0(CRC_OUT[12]),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .O(\TX_DATA_DEL14[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[13]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [13]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[13]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [13]));
  (* SOFT_HLUTNM = "soft_lutpair397" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[13]_i_2 
       (.I0(CRC_OUT[13]),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .O(\TX_DATA_DEL14[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[14]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [14]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[14]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[14]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [14]));
  (* SOFT_HLUTNM = "soft_lutpair396" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[14]_i_2 
       (.I0(CRC_OUT[14]),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .O(\TX_DATA_DEL14[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[15]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [15]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[15]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[15]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [15]));
  (* SOFT_HLUTNM = "soft_lutpair395" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[15]_i_3 
       (.I0(CRC_OUT[15]),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .O(\TX_DATA_DEL14[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hDFD0DFDFCFC0C0C0)) 
    \TX_DATA_DEL14[16]_i_1 
       (.I0(\TX_DATA_DEL14_reg[18] ),
        .I1(\TX_DATA_DEL14[16]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [16]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[16]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [16]));
  LUT6 #(
    .INIT(64'hB0F0B00000000000)) 
    \TX_DATA_DEL14[16]_i_2 
       (.I0(CRC_OUT[16]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[26] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00E2AAE2)) 
    \TX_DATA_DEL14[17]_i_1 
       (.I0(TX_DATA_DEL13[17]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[38] [17]),
        .I3(txstatplus_int0_out),
        .I4(\TX_DATA_DEL14_reg[18] ),
        .I5(\TX_DATA_DEL14[17]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [17]));
  LUT6 #(
    .INIT(64'hB0F0B00000000000)) 
    \TX_DATA_DEL14[17]_i_2 
       (.I0(CRC_OUT[17]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[21] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hE222FFFFE2220000)) 
    \TX_DATA_DEL14[18]_i_1 
       (.I0(TX_DATA_DEL13[18]),
        .I1(\TX_DATA_DEL14_reg[18] ),
        .I2(\TX_DATA_DEL14[18]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14[18]_i_3_n_0 ),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14_reg[18]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [18]));
  (* SOFT_HLUTNM = "soft_lutpair394" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \TX_DATA_DEL14[18]_i_2 
       (.I0(CRC_OUT[18]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[18]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair373" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \TX_DATA_DEL14[18]_i_3 
       (.I0(\TX_DATA_DEL14_reg[32] ),
        .I1(CRC_OUT[2]),
        .I2(fcs_enabled_int),
        .O(\TX_DATA_DEL14[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00E2AAE2)) 
    \TX_DATA_DEL14[19]_i_1 
       (.I0(TX_DATA_DEL13[19]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[38] [18]),
        .I3(txstatplus_int0_out),
        .I4(\TX_DATA_DEL14_reg[18] ),
        .I5(\TX_DATA_DEL14[19]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [19]));
  LUT6 #(
    .INIT(64'h8C0C800C00000000)) 
    \TX_DATA_DEL14[19]_i_2 
       (.I0(CRC_OUT[19]),
        .I1(\TX_DATA_DEL14_reg[21] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[3]),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[1]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [1]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[1]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [1]));
  (* SOFT_HLUTNM = "soft_lutpair395" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[1]_i_2 
       (.I0(CRC_OUT[1]),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .O(\TX_DATA_DEL14[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00E2AAE2)) 
    \TX_DATA_DEL14[20]_i_1 
       (.I0(TX_DATA_DEL13[20]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[38] [19]),
        .I3(txstatplus_int0_out),
        .I4(\TX_DATA_DEL14_reg[18] ),
        .I5(\TX_DATA_DEL14[20]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [20]));
  LUT6 #(
    .INIT(64'h8C0C800C00000000)) 
    \TX_DATA_DEL14[20]_i_2 
       (.I0(CRC_OUT[20]),
        .I1(\TX_DATA_DEL14_reg[21] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[4]),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00E2AAE2)) 
    \TX_DATA_DEL14[21]_i_1 
       (.I0(TX_DATA_DEL13[21]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[38] [20]),
        .I3(txstatplus_int0_out),
        .I4(\TX_DATA_DEL14_reg[18] ),
        .I5(\TX_DATA_DEL14[21]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [21]));
  LUT6 #(
    .INIT(64'h8C0C800C00000000)) 
    \TX_DATA_DEL14[21]_i_2 
       (.I0(CRC_OUT[21]),
        .I1(\TX_DATA_DEL14_reg[21] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[5]),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hDFD0DFDFCFC0C0C0)) 
    \TX_DATA_DEL14[22]_i_1 
       (.I0(\TX_DATA_DEL14_reg[18] ),
        .I1(\TX_DATA_DEL14[22]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [21]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[22]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [22]));
  LUT6 #(
    .INIT(64'h8C0C800C00000000)) 
    \TX_DATA_DEL14[22]_i_2 
       (.I0(CRC_OUT[22]),
        .I1(\TX_DATA_DEL14_reg[26] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[6]),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hDFD0DFDFCFC0C0C0)) 
    \TX_DATA_DEL14[23]_i_1 
       (.I0(\TX_DATA_DEL14_reg[18] ),
        .I1(\TX_DATA_DEL14[23]_i_3_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [22]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[23]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [23]));
  LUT6 #(
    .INIT(64'h8C0C800C00000000)) 
    \TX_DATA_DEL14[23]_i_3 
       (.I0(CRC_OUT[23]),
        .I1(\TX_DATA_DEL14_reg[26] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[7]),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \TX_DATA_DEL14[24]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[24]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [24]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[24]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [24]));
  LUT6 #(
    .INIT(64'hD1D1D1D1FCF030F0)) 
    \TX_DATA_DEL14[24]_i_2 
       (.I0(\TX_DATA_DEL14[24]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(TX_DATA_DEL13[24]),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFE00008002)) 
    \TX_DATA_DEL14[24]_i_3 
       (.I0(\TX_DATA_DEL14[56]_i_6_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(TX_DATA_VALID_DEL13__0[1]),
        .I3(TX_DATA_VALID_DEL13__0[0]),
        .I4(\TX_DATA_DEL14[57]_i_2_0 ),
        .I5(\TX_DATA_DEL14[8]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8FFFFBBB80000)) 
    \TX_DATA_DEL14[25]_i_1 
       (.I0(TX_DATA_DEL13[25]),
        .I1(TX_DATA_VALID_DEL13),
        .I2(\TX_DATA_DEL14[25]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14[25]_i_3_n_0 ),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14_reg[25] ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [25]));
  LUT5 #(
    .INIT(32'hC088C0C0)) 
    \TX_DATA_DEL14[25]_i_2 
       (.I0(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(TX_DATA_DEL13[25]),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1510555515100000)) 
    \TX_DATA_DEL14[25]_i_3 
       (.I0(\TX_DATA_DEL14_reg[58] ),
        .I1(\OVERFLOW_DATA[1]_i_3_n_0 ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(\TX_DATA_DEL14[9]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(TX_DATA_DEL13[25]),
        .O(\TX_DATA_DEL14[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFCACAFFFFFAFA)) 
    \TX_DATA_DEL14[26]_i_1 
       (.I0(append_end_frame),
        .I1(\TX_DATA_DEL14[26]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_VALID_DEL13),
        .I4(TX_DATA_DEL13[26]),
        .I5(\TX_DATA_DEL14[26]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [26]));
  LUT6 #(
    .INIT(64'h4000404040444040)) 
    \TX_DATA_DEL14[26]_i_2 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(TX_DATA_DEL13[26]),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[2]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FF00FFFFFF)) 
    \TX_DATA_DEL14[26]_i_3 
       (.I0(\OVERFLOW_DATA[2]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(\OVERFLOW_DATA[2]_i_3_n_0 ),
        .I3(\TX_DATA_DEL14_reg[26] ),
        .I4(TX_DATA_DEL13[26]),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \TX_DATA_DEL14[27]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[27]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [23]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[27]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [27]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \TX_DATA_DEL14[27]_i_2 
       (.I0(\TX_DATA_DEL14[27]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14[27]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[27]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFD01000101)) 
    \TX_DATA_DEL14[27]_i_3 
       (.I0(\TX_DATA_DEL14[3]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[57]_i_2_0 ),
        .I2(\TX_DATA_DEL14[57]_i_2_2 ),
        .I3(\TX_DATA_DEL14[57]_i_2_1 ),
        .I4(\TX_DATA_DEL14[63]_i_2_0 ),
        .I5(TX_DATA_DEL13[27]),
        .O(\TX_DATA_DEL14[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[27]_i_4 
       (.I0(\TX_DATA_DEL14[51]_i_6_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[27]),
        .O(\TX_DATA_DEL14[27]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[27]_i_5 
       (.I0(\TX_DATA_DEL14[11]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[27]),
        .O(\TX_DATA_DEL14[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \TX_DATA_DEL14[28]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[28]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [23]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[28]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [28]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \TX_DATA_DEL14[28]_i_2 
       (.I0(\TX_DATA_DEL14[28]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14[28]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[28]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFD01000101)) 
    \TX_DATA_DEL14[28]_i_3 
       (.I0(\TX_DATA_DEL14[4]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[57]_i_2_0 ),
        .I2(\TX_DATA_DEL14[57]_i_2_2 ),
        .I3(\TX_DATA_DEL14[57]_i_2_1 ),
        .I4(\TX_DATA_DEL14[63]_i_2_0 ),
        .I5(TX_DATA_DEL13[28]),
        .O(\TX_DATA_DEL14[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[28]_i_4 
       (.I0(\TX_DATA_DEL14[52]_i_5_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[28]),
        .O(\TX_DATA_DEL14[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[28]_i_5 
       (.I0(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[28]),
        .O(\TX_DATA_DEL14[28]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \TX_DATA_DEL14[29]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[29]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [23]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[29]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [29]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \TX_DATA_DEL14[29]_i_2 
       (.I0(\TX_DATA_DEL14[29]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14[29]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[29]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFD01000101)) 
    \TX_DATA_DEL14[29]_i_3 
       (.I0(\TX_DATA_DEL14[5]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[57]_i_2_0 ),
        .I2(\TX_DATA_DEL14[57]_i_2_2 ),
        .I3(\TX_DATA_DEL14[57]_i_2_1 ),
        .I4(\TX_DATA_DEL14[63]_i_2_0 ),
        .I5(TX_DATA_DEL13[29]),
        .O(\TX_DATA_DEL14[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[29]_i_4 
       (.I0(\TX_DATA_DEL14[53]_i_5_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[29]),
        .O(\TX_DATA_DEL14[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[29]_i_5 
       (.I0(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[29]),
        .O(\TX_DATA_DEL14[29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7F707F7F4F404040)) 
    \TX_DATA_DEL14[2]_i_1 
       (.I0(\TX_DATA_DEL14[2]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14_reg[0] ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [2]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[2]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [2]));
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[2]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[2]),
        .O(\TX_DATA_DEL14[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \TX_DATA_DEL14[30]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[30]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [23]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[30]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [30]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \TX_DATA_DEL14[30]_i_2 
       (.I0(\TX_DATA_DEL14[30]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14[30]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[30]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFD01000101)) 
    \TX_DATA_DEL14[30]_i_3 
       (.I0(\TX_DATA_DEL14[6]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[57]_i_2_0 ),
        .I2(\TX_DATA_DEL14[57]_i_2_2 ),
        .I3(\TX_DATA_DEL14[57]_i_2_1 ),
        .I4(\TX_DATA_DEL14[63]_i_2_0 ),
        .I5(TX_DATA_DEL13[30]),
        .O(\TX_DATA_DEL14[30]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[30]_i_4 
       (.I0(\TX_DATA_DEL14[54]_i_7_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[30]),
        .O(\TX_DATA_DEL14[30]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[30]_i_5 
       (.I0(\TX_DATA_DEL14[14]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[30]),
        .O(\TX_DATA_DEL14[30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \TX_DATA_DEL14[31]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[31]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [23]),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[31]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [31]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \TX_DATA_DEL14[31]_i_2 
       (.I0(\TX_DATA_DEL14[31]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14[31]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[31]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA20EF)) 
    \TX_DATA_DEL14[31]_i_3 
       (.I0(TX_DATA_DEL13[31]),
        .I1(\TX_DATA_DEL14[57]_i_2_1 ),
        .I2(\TX_DATA_DEL14[63]_i_2_0 ),
        .I3(\TX_DATA_DEL14[7]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14[57]_i_2_2 ),
        .I5(\TX_DATA_DEL14[57]_i_2_0 ),
        .O(\TX_DATA_DEL14[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[31]_i_4 
       (.I0(\TX_DATA_DEL14[55]_i_5_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[31]),
        .O(\TX_DATA_DEL14[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[31]_i_5 
       (.I0(\TX_DATA_DEL14[15]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(TX_DATA_DEL13[31]),
        .O(\TX_DATA_DEL14[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEFAFAA)) 
    \TX_DATA_DEL14[32]_i_1 
       (.I0(\TX_DATA_DEL14[32]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[32]),
        .I5(\TX_DATA_DEL14[32]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [32]));
  LUT6 #(
    .INIT(64'h20AA2AAA20002A00)) 
    \TX_DATA_DEL14[32]_i_2 
       (.I0(\TX_DATA_DEL14_reg[21] ),
        .I1(\OVERFLOW_DATA_reg[8] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\OVERFLOW_DATA[8]_i_3_n_0 ),
        .I5(TX_DATA_DEL13[32]),
        .O(\TX_DATA_DEL14[32]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC500C500FF000000)) 
    \TX_DATA_DEL14[32]_i_3 
       (.I0(\TX_DATA_DEL14[8]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14_reg[32]_0 ),
        .I4(TX_DATA_DEL13[32]),
        .I5(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[32]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8FFFFBBB80000)) 
    \TX_DATA_DEL14[33]_i_1 
       (.I0(TX_DATA_DEL13[33]),
        .I1(TX_DATA_VALID_DEL13),
        .I2(\TX_DATA_DEL14[33]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14[33]_i_3_n_0 ),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14_reg[33]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [33]));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \TX_DATA_DEL14[33]_i_2 
       (.I0(TX_DATA_DEL13[33]),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(\TX_DATA_DEL14[9]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[58] ),
        .O(\TX_DATA_DEL14[33]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0404045454540454)) 
    \TX_DATA_DEL14[33]_i_3 
       (.I0(\TX_DATA_DEL14_reg[58] ),
        .I1(TX_DATA_DEL13[33]),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14[33]_i_5_n_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14_reg[33] ),
        .O(\TX_DATA_DEL14[33]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair403" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[33]_i_5 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[17]),
        .O(\TX_DATA_DEL14[33]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEFEF4F40)) 
    \TX_DATA_DEL14[34]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[34]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[34]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [34]));
  LUT6 #(
    .INIT(64'h7C7F7F7F70734040)) 
    \TX_DATA_DEL14[34]_i_2 
       (.I0(\TX_DATA_DEL14[34]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(\TX_DATA_DEL14[50]_i_4_n_0 ),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(TX_DATA_DEL13[34]),
        .O(\TX_DATA_DEL14[34]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[34]_i_3 
       (.I0(\TX_DATA_DEL14[2]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\OVERFLOW_DATA[2]_i_3_n_0 ),
        .O(\TX_DATA_DEL14[34]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7770000)) 
    \TX_DATA_DEL14[35]_i_1 
       (.I0(\TX_DATA_DEL14[35]_i_2_n_0 ),
        .I1(txstatplus_int0_out),
        .I2(TX_DATA_VALID_DEL13),
        .I3(TX_DATA_DEL13[35]),
        .I4(\TX_DATA_DEL14_reg[39] ),
        .I5(\TX_DATA_DEL14[35]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [35]));
  LUT6 #(
    .INIT(64'h30703F7FFFFFFFFF)) 
    \TX_DATA_DEL14[35]_i_2 
       (.I0(CRC_OUT[19]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(TX_DATA_DEL13[35]),
        .I5(\TX_DATA_DEL14_reg[26] ),
        .O(\TX_DATA_DEL14[35]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC4C4C4FF80808080)) 
    \TX_DATA_DEL14[35]_i_3 
       (.I0(\TX_DATA_DEL14_reg[32] ),
        .I1(\TX_DATA_DEL14_reg[32]_0 ),
        .I2(\TX_DATA_DEL14[51]_i_4_n_0 ),
        .I3(append_end_frame),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[35]),
        .O(\TX_DATA_DEL14[35]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7770000)) 
    \TX_DATA_DEL14[36]_i_1 
       (.I0(\TX_DATA_DEL14[36]_i_2_n_0 ),
        .I1(txstatplus_int0_out),
        .I2(TX_DATA_VALID_DEL13),
        .I3(TX_DATA_DEL13[36]),
        .I4(\TX_DATA_DEL14_reg[39] ),
        .I5(\TX_DATA_DEL14[36]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [36]));
  LUT6 #(
    .INIT(64'h30703F7FFFFFFFFF)) 
    \TX_DATA_DEL14[36]_i_2 
       (.I0(CRC_OUT[20]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(TX_DATA_DEL13[36]),
        .I5(\TX_DATA_DEL14_reg[26] ),
        .O(\TX_DATA_DEL14[36]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC4C4C4FF80808080)) 
    \TX_DATA_DEL14[36]_i_3 
       (.I0(\TX_DATA_DEL14_reg[32] ),
        .I1(\TX_DATA_DEL14_reg[32]_0 ),
        .I2(\TX_DATA_DEL14[36]_i_4_n_0 ),
        .I3(append_end_frame),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[36]),
        .O(\TX_DATA_DEL14[36]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FF700004004)) 
    \TX_DATA_DEL14[36]_i_4 
       (.I0(\TX_DATA_DEL14[4]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[36]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7770000)) 
    \TX_DATA_DEL14[37]_i_1 
       (.I0(\TX_DATA_DEL14[37]_i_2_n_0 ),
        .I1(txstatplus_int0_out),
        .I2(TX_DATA_VALID_DEL13),
        .I3(TX_DATA_DEL13[37]),
        .I4(\TX_DATA_DEL14_reg[39] ),
        .I5(\TX_DATA_DEL14[37]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [37]));
  LUT6 #(
    .INIT(64'h30703F7FFFFFFFFF)) 
    \TX_DATA_DEL14[37]_i_2 
       (.I0(CRC_OUT[21]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(TX_DATA_DEL13[37]),
        .I5(\TX_DATA_DEL14_reg[26] ),
        .O(\TX_DATA_DEL14[37]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC4C4C4FF80808080)) 
    \TX_DATA_DEL14[37]_i_3 
       (.I0(\TX_DATA_DEL14_reg[32] ),
        .I1(\TX_DATA_DEL14_reg[32]_0 ),
        .I2(\TX_DATA_DEL14[37]_i_4_n_0 ),
        .I3(append_end_frame),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[37]),
        .O(\TX_DATA_DEL14[37]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FF700004004)) 
    \TX_DATA_DEL14[37]_i_4 
       (.I0(\TX_DATA_DEL14[5]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[37]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEF20000FEF2FEF2)) 
    \TX_DATA_DEL14[38]_i_1 
       (.I0(TX_DATA_DEL13[38]),
        .I1(append_end_frame),
        .I2(txstatplus_int0_out),
        .I3(\TX_DATA_DEL14_reg[38] [25]),
        .I4(\TX_DATA_DEL14[38]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14[38]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [38]));
  LUT6 #(
    .INIT(64'hFFFFA2FF00FF80FF)) 
    \TX_DATA_DEL14[38]_i_2 
       (.I0(\TX_DATA_DEL14_reg[58] ),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(\TX_DATA_DEL14[54]_i_4_n_0 ),
        .I3(txstatplus_int0_out),
        .I4(TX_DATA_VALID_DEL13),
        .I5(TX_DATA_DEL13[38]),
        .O(\TX_DATA_DEL14[38]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h30703F7FFFFFFFFF)) 
    \TX_DATA_DEL14[38]_i_3 
       (.I0(CRC_OUT[22]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(TX_DATA_DEL13[38]),
        .I5(\TX_DATA_DEL14_reg[26] ),
        .O(\TX_DATA_DEL14[38]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7770000)) 
    \TX_DATA_DEL14[39]_i_1 
       (.I0(\TX_DATA_DEL14[39]_i_2_n_0 ),
        .I1(txstatplus_int0_out),
        .I2(TX_DATA_VALID_DEL13),
        .I3(TX_DATA_DEL13[39]),
        .I4(\TX_DATA_DEL14_reg[39] ),
        .I5(\TX_DATA_DEL14[39]_i_4_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [39]));
  LUT6 #(
    .INIT(64'h303F707FFFFFFFFF)) 
    \TX_DATA_DEL14[39]_i_2 
       (.I0(CRC_OUT[23]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(TX_DATA_DEL13[39]),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14_reg[26] ),
        .O(\TX_DATA_DEL14[39]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC4C4C4FF80808080)) 
    \TX_DATA_DEL14[39]_i_4 
       (.I0(\TX_DATA_DEL14_reg[32] ),
        .I1(\TX_DATA_DEL14_reg[32]_0 ),
        .I2(\TX_DATA_DEL14[39]_i_6_n_0 ),
        .I3(append_end_frame),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[39]),
        .O(\TX_DATA_DEL14[39]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAA3A)) 
    \TX_DATA_DEL14[39]_i_6 
       (.I0(\TX_DATA_DEL14[15]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[7]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[63]_i_2_0 ),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .I5(TX_DATA_VALID_DEL13__0[5]),
        .O(\TX_DATA_DEL14[39]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB0F008888)) 
    \TX_DATA_DEL14[3]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [3]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14[3]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[0] ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[3]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [3]));
  (* SOFT_HLUTNM = "soft_lutpair391" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[3]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[3]),
        .O(\TX_DATA_DEL14[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFF54FF5400)) 
    \TX_DATA_DEL14[40]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[40]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[40]_i_3_n_0 ),
        .I3(txstatplus_int0_out),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[40]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [40]));
  LUT6 #(
    .INIT(64'h0000A808AAAAA808)) 
    \TX_DATA_DEL14[40]_i_2 
       (.I0(\TX_DATA_DEL14_reg[58] ),
        .I1(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(TX_DATA_DEL13[40]),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[56]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[40]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000FBFB0000FF00)) 
    \TX_DATA_DEL14[40]_i_3 
       (.I0(CRC_OUT[24]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(TX_DATA_DEL13[40]),
        .I4(\TX_DATA_DEL14_reg[58] ),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[40]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEFEF4F40)) 
    \TX_DATA_DEL14[41]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[41]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[41]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [41]));
  LUT6 #(
    .INIT(64'hB8FFB800B8FFB8FF)) 
    \TX_DATA_DEL14[41]_i_2 
       (.I0(\TX_DATA_DEL14[57]_i_4_n_0 ),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(\TX_DATA_DEL14[41]_i_3_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58] ),
        .I4(\TX_DATA_DEL14[41]_i_4_n_0 ),
        .I5(\TX_DATA_DEL14_reg[41] ),
        .O(\TX_DATA_DEL14[41]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[41]_i_3 
       (.I0(TX_DATA_DEL13[41]),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[41]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000FD0000)) 
    \TX_DATA_DEL14[41]_i_4 
       (.I0(\OVERFLOW_DATA_reg[8] ),
        .I1(\TX_DATA_DEL14[57]_i_2_2 ),
        .I2(\TX_DATA_DEL14[57]_i_2_0 ),
        .I3(\TX_DATA_DEL14[57]_i_2_1 ),
        .I4(\TX_DATA_DEL14[63]_i_2_0 ),
        .I5(\OVERFLOW_DATA[1]_i_3_n_0 ),
        .O(\TX_DATA_DEL14[41]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFF54FF5400)) 
    \TX_DATA_DEL14[42]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[42]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[42]_i_3_n_0 ),
        .I3(txstatplus_int0_out),
        .I4(append_end_frame),
        .I5(TX_DATA_DEL13[42]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [42]));
  LUT6 #(
    .INIT(64'h0000A202AAAAA202)) 
    \TX_DATA_DEL14[42]_i_2 
       (.I0(\TX_DATA_DEL14_reg[58] ),
        .I1(\TX_DATA_DEL14[2]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(TX_DATA_DEL13[42]),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[42]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[42]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000FBFB0000FF00)) 
    \TX_DATA_DEL14[42]_i_3 
       (.I0(CRC_OUT[26]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(TX_DATA_DEL13[42]),
        .I4(\TX_DATA_DEL14_reg[58] ),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[42]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[42]_i_4 
       (.I0(\OVERFLOW_DATA[2]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[50]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[42]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF44444444)) 
    \TX_DATA_DEL14[43]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[43]),
        .I2(\TX_DATA_DEL14[43]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58] ),
        .I4(\TX_DATA_DEL14[43]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14_reg[58]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [43]));
  LUT6 #(
    .INIT(64'h0F000FFF55CC55CC)) 
    \TX_DATA_DEL14[43]_i_2 
       (.I0(TX_DATA_DEL13[43]),
        .I1(\TX_DATA_DEL14[3]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[11]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14[43]_i_4_n_0 ),
        .I5(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[43]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4F7F00004F7FFFFF)) 
    \TX_DATA_DEL14[43]_i_3 
       (.I0(txstatplus_int),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[27]),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(TX_DATA_DEL13[43]),
        .O(\TX_DATA_DEL14[43]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair378" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[43]_i_4 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[19]),
        .O(\TX_DATA_DEL14[43]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF44444444)) 
    \TX_DATA_DEL14[44]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[44]),
        .I2(\TX_DATA_DEL14[44]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58] ),
        .I4(\TX_DATA_DEL14[44]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14_reg[58]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [44]));
  LUT6 #(
    .INIT(64'h0F000FFF55CC55CC)) 
    \TX_DATA_DEL14[44]_i_2 
       (.I0(TX_DATA_DEL13[44]),
        .I1(\TX_DATA_DEL14[4]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14[52]_i_4_n_0 ),
        .I5(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[44]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4F7F00004F7FFFFF)) 
    \TX_DATA_DEL14[44]_i_3 
       (.I0(txstatplus_int),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[28]),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(TX_DATA_DEL13[44]),
        .O(\TX_DATA_DEL14[44]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF44444444)) 
    \TX_DATA_DEL14[45]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[45]),
        .I2(\TX_DATA_DEL14[45]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58] ),
        .I4(\TX_DATA_DEL14[45]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14_reg[58]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [45]));
  LUT6 #(
    .INIT(64'h0F000FFF55CC55CC)) 
    \TX_DATA_DEL14[45]_i_2 
       (.I0(TX_DATA_DEL13[45]),
        .I1(\TX_DATA_DEL14[5]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14[53]_i_4_n_0 ),
        .I5(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[45]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4F7F00004F7FFFFF)) 
    \TX_DATA_DEL14[45]_i_3 
       (.I0(txstatplus_int),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[29]),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(TX_DATA_DEL13[45]),
        .O(\TX_DATA_DEL14[45]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF44444444)) 
    \TX_DATA_DEL14[46]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[46]),
        .I2(\TX_DATA_DEL14[46]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58] ),
        .I4(\TX_DATA_DEL14[46]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14_reg[58]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [46]));
  LUT6 #(
    .INIT(64'h553355330FFF0F00)) 
    \TX_DATA_DEL14[46]_i_2 
       (.I0(\TX_DATA_DEL14[14]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[46]_i_4_n_0 ),
        .I2(TX_DATA_DEL13[46]),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\TX_DATA_DEL14[6]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[46]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4F7F00004F7FFFFF)) 
    \TX_DATA_DEL14[46]_i_3 
       (.I0(txstatplus_int),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(fcs_enabled_int),
        .I3(CRC_OUT[30]),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(TX_DATA_DEL13[46]),
        .O(\TX_DATA_DEL14[46]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair375" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[46]_i_4 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[22]),
        .O(\TX_DATA_DEL14[46]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F0F44444444)) 
    \TX_DATA_DEL14[47]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[47]),
        .I2(\TX_DATA_DEL14[47]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[47] ),
        .I4(\TX_DATA_DEL14[47]_i_4_n_0 ),
        .I5(\TX_DATA_DEL14_reg[58]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [47]));
  LUT6 #(
    .INIT(64'h00002A20AAAA2A20)) 
    \TX_DATA_DEL14[47]_i_2 
       (.I0(\TX_DATA_DEL14_reg[58] ),
        .I1(TX_DATA_DEL13[47]),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(\TX_DATA_DEL14[7]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[63]_i_6_n_0 ),
        .O(\TX_DATA_DEL14[47]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair383" *) 
  LUT5 #(
    .INIT(32'h4FFF7FFF)) 
    \TX_DATA_DEL14[47]_i_4 
       (.I0(txstatplus_int),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(\TX_DATA_DEL14_reg[50] ),
        .I3(fcs_enabled_int),
        .I4(CRC_OUT[31]),
        .O(\TX_DATA_DEL14[47]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEFEF4F40)) 
    \TX_DATA_DEL14[48]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[48]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[48]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [48]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \TX_DATA_DEL14[48]_i_2 
       (.I0(\TX_DATA_DEL14[48]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[48]_i_4_n_0 ),
        .I2(\TX_DATA_DEL14_reg[58] ),
        .I3(\TX_DATA_DEL14_reg[48] ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14_reg[48]_0 ),
        .O(\TX_DATA_DEL14[48]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h5555555535555535)) 
    \TX_DATA_DEL14[48]_i_3 
       (.I0(\TX_DATA_DEL14[56]_i_6_n_0 ),
        .I1(\OVERFLOW_DATA[8]_i_3_n_0 ),
        .I2(\TX_DATA_DEL14[63]_i_2_0 ),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .I5(TX_DATA_VALID_DEL13__0[5]),
        .O(\TX_DATA_DEL14[48]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h55555555C55555C5)) 
    \TX_DATA_DEL14[48]_i_4 
       (.I0(\TX_DATA_DEL14[8]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[63]_i_2_0 ),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .I5(TX_DATA_VALID_DEL13__0[5]),
        .O(\TX_DATA_DEL14[48]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEFEF4F40)) 
    \TX_DATA_DEL14[49]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[49]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[49]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [49]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \TX_DATA_DEL14[49]_i_2 
       (.I0(\TX_DATA_DEL14[49]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[49]_i_4_n_0 ),
        .I2(\TX_DATA_DEL14_reg[58] ),
        .I3(\TX_DATA_DEL14_reg[49] ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14_reg[49]_0 ),
        .O(\TX_DATA_DEL14[49]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h555515515555D55D)) 
    \TX_DATA_DEL14[49]_i_3 
       (.I0(\OVERFLOW_DATA[1]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[33]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[49]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[49]_i_4 
       (.I0(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[9]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[49]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB0F008888)) 
    \TX_DATA_DEL14[4]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [4]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14[4]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[0] ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[4]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [4]));
  (* SOFT_HLUTNM = "soft_lutpair407" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[4]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[4]),
        .O(\TX_DATA_DEL14[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hCFCFCFC0FFAAFFAA)) 
    \TX_DATA_DEL14[50]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(\TX_DATA_DEL14[50]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14_reg[58] ),
        .I3(TX_DATA_DEL13[50]),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(\TX_DATA_DEL14_reg[58]_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [50]));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \TX_DATA_DEL14[50]_i_2 
       (.I0(\TX_DATA_DEL14[50]_i_4_n_0 ),
        .I1(\OVERFLOW_DATA[2]_i_2_n_0 ),
        .I2(\TX_DATA_DEL14[2]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[50] ),
        .I4(\OVERFLOW_DATA[2]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14_reg[32] ),
        .O(\TX_DATA_DEL14[50]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair394" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[50]_i_4 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[18]),
        .O(\TX_DATA_DEL14[50]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE040EF40)) 
    \TX_DATA_DEL14[51]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[51]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[51]),
        .I4(append_end_frame),
        .O(\TX_DATA_VALID_DEL13_reg[7] [51]));
  LUT6 #(
    .INIT(64'hAFAFCFCFA0A0C0CF)) 
    \TX_DATA_DEL14[51]_i_2 
       (.I0(\TX_DATA_DEL14[51]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[51]_i_4_n_0 ),
        .I2(\TX_DATA_DEL14_reg[58] ),
        .I3(\TX_DATA_DEL14_reg[54] ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14_reg[51] ),
        .O(\TX_DATA_DEL14[51]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[51]_i_3 
       (.I0(\TX_DATA_DEL14[43]_i_4_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[51]_i_6_n_0 ),
        .O(\TX_DATA_DEL14[51]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FF700004004)) 
    \TX_DATA_DEL14[51]_i_4 
       (.I0(\TX_DATA_DEL14[3]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[11]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[51]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair402" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[51]_i_6 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[27]),
        .O(\TX_DATA_DEL14[51]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF404F4F4F4040404)) 
    \TX_DATA_DEL14[52]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[52]),
        .I2(\TX_DATA_DEL14_reg[58]_0 ),
        .I3(\TX_DATA_DEL14[52]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[58] ),
        .I5(\TX_DATA_DEL14_reg[52] ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [52]));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \TX_DATA_DEL14[52]_i_2 
       (.I0(\TX_DATA_DEL14[52]_i_4_n_0 ),
        .I1(\TX_DATA_DEL14[52]_i_5_n_0 ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(\TX_DATA_DEL14[4]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[52]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair381" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[52]_i_4 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[20]),
        .O(\TX_DATA_DEL14[52]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair401" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[52]_i_5 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[28]),
        .O(\TX_DATA_DEL14[52]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF404F4F4F4040404)) 
    \TX_DATA_DEL14[53]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[53]),
        .I2(\TX_DATA_DEL14_reg[58]_0 ),
        .I3(\TX_DATA_DEL14[53]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[58] ),
        .I5(\TX_DATA_DEL14_reg[53] ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [53]));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \TX_DATA_DEL14[53]_i_2 
       (.I0(\TX_DATA_DEL14[53]_i_4_n_0 ),
        .I1(\TX_DATA_DEL14[53]_i_5_n_0 ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(\TX_DATA_DEL14[5]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .I5(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[53]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair374" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[53]_i_4 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[21]),
        .O(\TX_DATA_DEL14[53]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair399" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[53]_i_5 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[29]),
        .O(\TX_DATA_DEL14[53]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE040EF40)) 
    \TX_DATA_DEL14[54]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[54]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[54]),
        .I4(append_end_frame),
        .O(\TX_DATA_VALID_DEL13_reg[7] [54]));
  LUT6 #(
    .INIT(64'hAFAFCFCFA0A0C0CF)) 
    \TX_DATA_DEL14[54]_i_2 
       (.I0(\TX_DATA_DEL14[54]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[54]_i_4_n_0 ),
        .I2(\TX_DATA_DEL14_reg[58] ),
        .I3(\TX_DATA_DEL14_reg[54] ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14_reg[54]_0 ),
        .O(\TX_DATA_DEL14[54]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEAAEAAAA2AA2)) 
    \TX_DATA_DEL14[54]_i_3 
       (.I0(\TX_DATA_DEL14[54]_i_7_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[46]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[54]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FF700004004)) 
    \TX_DATA_DEL14[54]_i_4 
       (.I0(\TX_DATA_DEL14[6]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[14]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[54]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair401" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[54]_i_7 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[30]),
        .O(\TX_DATA_DEL14[54]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF404F4F4F4040404)) 
    \TX_DATA_DEL14[55]_i_1 
       (.I0(\TX_DATA_DEL14_reg[58]_1 ),
        .I1(TX_DATA_DEL13[55]),
        .I2(\TX_DATA_DEL14_reg[58]_0 ),
        .I3(\TX_DATA_DEL14[55]_i_2_n_0 ),
        .I4(\TX_DATA_DEL14_reg[58] ),
        .I5(\TX_DATA_DEL14_reg[55] ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [55]));
  LUT6 #(
    .INIT(64'hA0A0AFAFCFC0CFC0)) 
    \TX_DATA_DEL14[55]_i_2 
       (.I0(\TX_DATA_DEL14[55]_i_4_n_0 ),
        .I1(\TX_DATA_DEL14[55]_i_5_n_0 ),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(\TX_DATA_DEL14[15]_i_3_n_0 ),
        .I4(\TX_DATA_DEL14[7]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[55]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair377" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[55]_i_4 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[23]),
        .O(\TX_DATA_DEL14[55]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair383" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[55]_i_5 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[31]),
        .O(\TX_DATA_DEL14[55]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFCFC0)) 
    \TX_DATA_DEL14[56]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[56]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[56]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [56]));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \TX_DATA_DEL14[56]_i_2 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[56]_i_3_n_0 ),
        .I2(\TX_DATA_DEL14_reg[58] ),
        .I3(\TX_DATA_DEL14[56]_i_4_n_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[56]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[56]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h3335333500003335)) 
    \TX_DATA_DEL14[56]_i_3 
       (.I0(\TX_DATA_DEL14[0]_i_2_n_0 ),
        .I1(TX_DATA_DEL13[56]),
        .I2(\TX_DATA_DEL14[57]_i_2_0 ),
        .I3(\TX_DATA_DEL14[57]_i_2_2 ),
        .I4(\TX_DATA_DEL14[63]_i_2_0 ),
        .I5(\TX_DATA_DEL14[57]_i_2_1 ),
        .O(\TX_DATA_DEL14[56]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[56]_i_4 
       (.I0(\TX_DATA_DEL14[8]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\OVERFLOW_DATA[8]_i_3_n_0 ),
        .O(\TX_DATA_DEL14[56]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[56]_i_5 
       (.I0(\TX_DATA_DEL14[56]_i_6_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\OVERFLOW_DATA_reg[8] ),
        .O(\TX_DATA_DEL14[56]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair386" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[56]_i_6 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[24]),
        .O(\TX_DATA_DEL14[56]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEFEF4F40)) 
    \TX_DATA_DEL14[57]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[57]_i_2_n_0 ),
        .I2(txstatplus_int0_out),
        .I3(append_end_frame),
        .I4(TX_DATA_DEL13[57]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [57]));
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \TX_DATA_DEL14[57]_i_2 
       (.I0(\TX_DATA_DEL14[57]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14_reg[32] ),
        .I2(\TX_DATA_DEL14[57]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58] ),
        .I4(\TX_DATA_DEL14[57]_i_5_n_0 ),
        .I5(\TX_DATA_DEL14_reg[57] ),
        .O(\TX_DATA_DEL14[57]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00004004FFFF7FF7)) 
    \TX_DATA_DEL14[57]_i_3 
       (.I0(\OVERFLOW_DATA[1]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14_reg[33] ),
        .O(\TX_DATA_DEL14[57]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5555D55D55551551)) 
    \TX_DATA_DEL14[57]_i_4 
       (.I0(\TX_DATA_DEL14[33]_i_5_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[9]_i_2_n_0 ),
        .O(\TX_DATA_DEL14[57]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \TX_DATA_DEL14[57]_i_5 
       (.I0(\TX_DATA_DEL14[1]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(\TX_DATA_DEL14[57]_i_2_1 ),
        .I3(\TX_DATA_DEL14[57]_i_2_2 ),
        .I4(\TX_DATA_DEL14[57]_i_2_0 ),
        .O(\TX_DATA_DEL14[57]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \TX_DATA_DEL14[58]_i_1 
       (.I0(\TX_DATA_DEL14[58]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14_reg[58] ),
        .I2(\TX_DATA_DEL14[58]_i_4_n_0 ),
        .I3(\TX_DATA_DEL14_reg[58]_0 ),
        .I4(TX_DATA_DEL13[58]),
        .I5(\TX_DATA_DEL14_reg[58]_1 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [58]));
  LUT6 #(
    .INIT(64'hFA0AFFFFFCFCFFFF)) 
    \TX_DATA_DEL14[58]_i_2 
       (.I0(CRC_OUT[10]),
        .I1(CRC_OUT[18]),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(CRC_OUT[26]),
        .I4(fcs_enabled_int),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[58]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair373" *) 
  LUT5 #(
    .INIT(32'hFFFFBFB0)) 
    \TX_DATA_DEL14[58]_i_4 
       (.I0(CRC_OUT[2]),
        .I1(fcs_enabled_int),
        .I2(\TX_DATA_DEL14_reg[32] ),
        .I3(TX_DATA_DEL13[58]),
        .I4(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[58]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEFAA)) 
    \TX_DATA_DEL14[59]_i_1 
       (.I0(\TX_DATA_DEL14[59]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[59]),
        .I4(append_end_frame),
        .I5(\TX_DATA_DEL14[59]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [59]));
  LUT6 #(
    .INIT(64'hC400FF00C4000000)) 
    \TX_DATA_DEL14[59]_i_2 
       (.I0(\TX_DATA_DEL14_reg[50] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[27]),
        .I3(\TX_DATA_DEL14_reg[32]_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[59]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[59]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00E233E200000000)) 
    \TX_DATA_DEL14[59]_i_3 
       (.I0(TX_DATA_DEL13[59]),
        .I1(\TX_DATA_DEL14_reg[50] ),
        .I2(\OVERFLOW_DATA_reg[8] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[3]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[21] ),
        .O(\TX_DATA_DEL14[59]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[59]_i_4 
       (.I0(\TX_DATA_DEL14[11]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[43]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[59]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB0F008888)) 
    \TX_DATA_DEL14[5]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [5]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14[5]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[0] ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[5]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [5]));
  (* SOFT_HLUTNM = "soft_lutpair407" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[5]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[5]),
        .O(\TX_DATA_DEL14[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEFAA)) 
    \TX_DATA_DEL14[60]_i_1 
       (.I0(\TX_DATA_DEL14[60]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[60]),
        .I4(append_end_frame),
        .I5(\TX_DATA_DEL14[60]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [60]));
  LUT6 #(
    .INIT(64'hC400FF00C4000000)) 
    \TX_DATA_DEL14[60]_i_2 
       (.I0(\TX_DATA_DEL14_reg[50] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[28]),
        .I3(\TX_DATA_DEL14_reg[32]_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[60]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[60]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00E233E200000000)) 
    \TX_DATA_DEL14[60]_i_3 
       (.I0(TX_DATA_DEL13[60]),
        .I1(\TX_DATA_DEL14_reg[50] ),
        .I2(\OVERFLOW_DATA_reg[8] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[4]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[21] ),
        .O(\TX_DATA_DEL14[60]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[60]_i_4 
       (.I0(\TX_DATA_DEL14[12]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[52]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[60]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEFAA)) 
    \TX_DATA_DEL14[61]_i_1 
       (.I0(\TX_DATA_DEL14[61]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[61]),
        .I4(append_end_frame),
        .I5(\TX_DATA_DEL14[61]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [61]));
  LUT6 #(
    .INIT(64'hC0880088CC880088)) 
    \TX_DATA_DEL14[61]_i_2 
       (.I0(\TX_DATA_DEL14[61]_i_4_n_0 ),
        .I1(\TX_DATA_DEL14_reg[32]_0 ),
        .I2(CRC_OUT[29]),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(fcs_enabled_int),
        .I5(\TX_DATA_DEL14_reg[50] ),
        .O(\TX_DATA_DEL14[61]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00E233E200000000)) 
    \TX_DATA_DEL14[61]_i_3 
       (.I0(TX_DATA_DEL13[61]),
        .I1(\TX_DATA_DEL14_reg[50] ),
        .I2(\OVERFLOW_DATA_reg[8] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[5]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[21] ),
        .O(\TX_DATA_DEL14[61]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[61]_i_4 
       (.I0(\TX_DATA_DEL14[13]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[53]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[61]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEFAA)) 
    \TX_DATA_DEL14[62]_i_1 
       (.I0(\TX_DATA_DEL14[62]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[62]),
        .I4(append_end_frame),
        .I5(\TX_DATA_DEL14[62]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [62]));
  LUT6 #(
    .INIT(64'h00E233E200000000)) 
    \TX_DATA_DEL14[62]_i_2 
       (.I0(TX_DATA_DEL13[62]),
        .I1(\TX_DATA_DEL14_reg[50] ),
        .I2(\OVERFLOW_DATA_reg[8] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[6]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[21] ),
        .O(\TX_DATA_DEL14[62]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC400FF00C4000000)) 
    \TX_DATA_DEL14[62]_i_3 
       (.I0(\TX_DATA_DEL14_reg[50] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[30]),
        .I3(\TX_DATA_DEL14_reg[32]_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[62]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[62]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[62]_i_4 
       (.I0(\TX_DATA_DEL14[14]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[46]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[62]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEFAA)) 
    \TX_DATA_DEL14[63]_i_1 
       (.I0(\TX_DATA_DEL14[63]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(txstatplus_int0_out),
        .I3(TX_DATA_DEL13[63]),
        .I4(append_end_frame),
        .I5(\TX_DATA_DEL14[63]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [63]));
  LUT6 #(
    .INIT(64'hC400FF00C4000000)) 
    \TX_DATA_DEL14[63]_i_2 
       (.I0(\TX_DATA_DEL14_reg[50] ),
        .I1(fcs_enabled_int),
        .I2(CRC_OUT[31]),
        .I3(\TX_DATA_DEL14_reg[32]_0 ),
        .I4(\TX_DATA_DEL14_reg[32] ),
        .I5(\TX_DATA_DEL14[63]_i_6_n_0 ),
        .O(\TX_DATA_DEL14[63]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00E233E200000000)) 
    \TX_DATA_DEL14[63]_i_3 
       (.I0(TX_DATA_DEL13[63]),
        .I1(\TX_DATA_DEL14_reg[50] ),
        .I2(\OVERFLOW_DATA_reg[8] ),
        .I3(\TX_DATA_DEL14_reg[32] ),
        .I4(\TX_DATA_DEL14[7]_i_2_n_0 ),
        .I5(\TX_DATA_DEL14_reg[21] ),
        .O(\TX_DATA_DEL14[63]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFB00008008)) 
    \TX_DATA_DEL14[63]_i_6 
       (.I0(\TX_DATA_DEL14[15]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_2_0 ),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .I5(\TX_DATA_DEL14[55]_i_4_n_0 ),
        .O(\TX_DATA_DEL14[63]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB0F008888)) 
    \TX_DATA_DEL14[6]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [6]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14[6]_i_2_n_0 ),
        .I3(\TX_DATA_DEL14_reg[0] ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[6]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [6]));
  (* SOFT_HLUTNM = "soft_lutpair406" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[6]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[6]),
        .O(\TX_DATA_DEL14[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB00F08888)) 
    \TX_DATA_DEL14[7]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [7]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(\TX_DATA_DEL14[7]_i_2_n_0 ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[7]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [7]));
  (* SOFT_HLUTNM = "soft_lutpair406" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[7]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[7]),
        .O(\TX_DATA_DEL14[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFBBBB00F08888)) 
    \TX_DATA_DEL14[8]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [8]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(\TX_DATA_DEL14[8]_i_2_n_0 ),
        .I4(txstatplus_int0_out),
        .I5(TX_DATA_DEL13[8]),
        .O(\TX_DATA_VALID_DEL13_reg[7] [8]));
  (* SOFT_HLUTNM = "soft_lutpair405" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[8]_i_2 
       (.I0(fcs_enabled_int),
        .I1(CRC_OUT[8]),
        .O(\TX_DATA_DEL14[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0BB880F00BB88)) 
    \TX_DATA_DEL14[9]_i_1 
       (.I0(\TX_DATA_DEL14_reg[38] [9]),
        .I1(append_end_frame),
        .I2(\TX_DATA_DEL14_reg[0] ),
        .I3(TX_DATA_DEL13[9]),
        .I4(txstatplus_int0_out),
        .I5(\TX_DATA_DEL14[9]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL13_reg[7] [9]));
  (* SOFT_HLUTNM = "soft_lutpair396" *) 
  LUT3 #(
    .INIT(8'hC5)) 
    \TX_DATA_DEL14[9]_i_2 
       (.I0(txstatplus_int),
        .I1(CRC_OUT[9]),
        .I2(fcs_enabled_int),
        .O(\TX_DATA_DEL14[9]_i_2_n_0 ));
endmodule

(* ORIG_REF_NAME = "CRC32_D8" *) 
module switch_elements_CRC32_D8_4
   (small_error_reg,
    D,
    small_error,
    large_error,
    Q,
    do_crc_check,
    wait_crc_check,
    \CRC_OUT_reg[30]_0 ,
    \CRC_OUT_reg[19]_0 ,
    \CRC_OUT_reg[31]_0 ,
    clk_i,
    reset_dcm);
  output small_error_reg;
  output [0:0]D;
  input small_error;
  input large_error;
  input [0:0]Q;
  input do_crc_check;
  input wait_crc_check;
  input [7:0]\CRC_OUT_reg[30]_0 ;
  input \CRC_OUT_reg[19]_0 ;
  input [31:0]\CRC_OUT_reg[31]_0 ;
  input clk_i;
  input reset_dcm;

  wire \CRC_OUT[10]_i_2__0_n_0 ;
  wire \CRC_OUT[10]_i_3__0_n_0 ;
  wire \CRC_OUT[11]_i_2__0_n_0 ;
  wire \CRC_OUT[12]_i_2__0_n_0 ;
  wire \CRC_OUT[13]_i_2__0_n_0 ;
  wire \CRC_OUT[13]_i_3__0_n_0 ;
  wire \CRC_OUT[13]_i_4__1_n_0 ;
  wire \CRC_OUT[14]_i_2__2_n_0 ;
  wire \CRC_OUT[14]_i_3__0_n_0 ;
  wire \CRC_OUT[15]_i_2__0_n_0 ;
  wire \CRC_OUT[15]_i_3__0_n_0 ;
  wire \CRC_OUT[16]_i_2__0_n_0 ;
  wire \CRC_OUT[16]_i_3__0_n_0 ;
  wire \CRC_OUT[16]_i_4__0_n_0 ;
  wire \CRC_OUT[17]_i_2__0_n_0 ;
  wire \CRC_OUT[18]_i_2__1_n_0 ;
  wire \CRC_OUT[18]_i_3__0_n_0 ;
  wire \CRC_OUT[19]_i_2__0_n_0 ;
  wire \CRC_OUT[23]_i_2__0_n_0 ;
  wire \CRC_OUT[24]_i_2__0_n_0 ;
  wire \CRC_OUT[24]_i_3__0_n_0 ;
  wire \CRC_OUT[24]_i_4__0_n_0 ;
  wire \CRC_OUT[25]_i_2__0_n_0 ;
  wire \CRC_OUT[26]_i_2__0_n_0 ;
  wire \CRC_OUT[27]_i_2__0_n_0 ;
  wire \CRC_OUT[28]_i_2__0_n_0 ;
  wire \CRC_OUT[29]_i_2__0_n_0 ;
  wire \CRC_OUT[2]_i_2__0_n_0 ;
  wire \CRC_OUT[30]_i_2__0_n_0 ;
  wire \CRC_OUT[3]_i_2__2_n_0 ;
  wire \CRC_OUT[4]_i_2__0_n_0 ;
  wire \CRC_OUT[5]_i_2__0_n_0 ;
  wire \CRC_OUT[5]_i_3__1_n_0 ;
  wire \CRC_OUT[6]_i_2__0_n_0 ;
  wire \CRC_OUT[7]_i_2__0_n_0 ;
  wire \CRC_OUT[9]_i_2__0_n_0 ;
  wire \CRC_OUT_reg[19]_0 ;
  wire [7:0]\CRC_OUT_reg[30]_0 ;
  wire [31:0]\CRC_OUT_reg[31]_0 ;
  wire [0:0]D;
  wire [0:0]Q;
  wire clk_i;
  wire [31:0]crc_from_8;
  wire do_crc_check;
  wire good_frame_get_i_3_n_0;
  wire large_error;
  wire [31:0]p_1_in;
  wire reset_dcm;
  wire \rxStatRegPlus[1]_i_10_n_0 ;
  wire \rxStatRegPlus[1]_i_2_n_0 ;
  wire \rxStatRegPlus[1]_i_3_n_0 ;
  wire \rxStatRegPlus[1]_i_4_n_0 ;
  wire \rxStatRegPlus[1]_i_5_n_0 ;
  wire \rxStatRegPlus[1]_i_6_n_0 ;
  wire \rxStatRegPlus[1]_i_7_n_0 ;
  wire \rxStatRegPlus[1]_i_8_n_0 ;
  wire \rxStatRegPlus[1]_i_9_n_0 ;
  wire small_error;
  wire small_error_reg;
  wire wait_crc_check;

  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[0]_i_1__0 
       (.I0(crc_from_8[24]),
        .I1(\CRC_OUT_reg[30]_0 [0]),
        .I2(crc_from_8[30]),
        .I3(\CRC_OUT_reg[30]_0 [6]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [0]),
        .O(p_1_in[0]));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[10]_i_1__0 
       (.I0(\CRC_OUT[10]_i_2__0_n_0 ),
        .I1(\CRC_OUT_reg[30]_0 [5]),
        .I2(crc_from_8[29]),
        .I3(\CRC_OUT[10]_i_3__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [10]),
        .O(p_1_in[10]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[10]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[24]),
        .I2(\CRC_OUT_reg[30]_0 [0]),
        .O(\CRC_OUT[10]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[10]_i_3__0 
       (.I0(crc_from_8[26]),
        .I1(\CRC_OUT_reg[30]_0 [3]),
        .I2(crc_from_8[2]),
        .I3(crc_from_8[27]),
        .O(\CRC_OUT[10]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[11]_i_1__0 
       (.I0(crc_from_8[3]),
        .I1(\CRC_OUT[11]_i_2__0_n_0 ),
        .I2(\CRC_OUT_reg[30]_0 [3]),
        .I3(\CRC_OUT_reg[30]_0 [4]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [11]),
        .O(p_1_in[11]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_2__0 
       (.I0(crc_from_8[27]),
        .I1(crc_from_8[28]),
        .I2(\CRC_OUT_reg[30]_0 [0]),
        .I3(crc_from_8[24]),
        .I4(crc_from_8[25]),
        .I5(\CRC_OUT_reg[30]_0 [1]),
        .O(\CRC_OUT[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[12]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [4]),
        .I1(\CRC_OUT[23]_i_2__0_n_0 ),
        .I2(\CRC_OUT[14]_i_2__2_n_0 ),
        .I3(\CRC_OUT[12]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [12]),
        .O(p_1_in[12]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[12]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [5]),
        .I1(\CRC_OUT_reg[30]_0 [6]),
        .I2(crc_from_8[29]),
        .I3(crc_from_8[28]),
        .I4(crc_from_8[4]),
        .O(\CRC_OUT[12]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[13]_i_1__0 
       (.I0(\CRC_OUT[13]_i_2__0_n_0 ),
        .I1(\CRC_OUT_reg[30]_0 [5]),
        .I2(\CRC_OUT[13]_i_3__0_n_0 ),
        .I3(\CRC_OUT[13]_i_4__1_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [13]),
        .O(p_1_in[13]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[5]),
        .I2(\CRC_OUT[24]_i_4__0_n_0 ),
        .I3(crc_from_8[26]),
        .I4(crc_from_8[27]),
        .I5(\CRC_OUT_reg[30]_0 [3]),
        .O(\CRC_OUT[13]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[13]_i_3__0 
       (.I0(\CRC_OUT_reg[30]_0 [7]),
        .I1(\CRC_OUT_reg[30]_0 [6]),
        .O(\CRC_OUT[13]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \CRC_OUT[13]_i_4__1 
       (.I0(crc_from_8[30]),
        .I1(crc_from_8[31]),
        .I2(crc_from_8[29]),
        .O(\CRC_OUT[13]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[14]_i_1__0 
       (.I0(crc_from_8[31]),
        .I1(\CRC_OUT[30]_i_2__0_n_0 ),
        .I2(\CRC_OUT[14]_i_2__2_n_0 ),
        .I3(\CRC_OUT[14]_i_3__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [14]),
        .O(p_1_in[14]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \CRC_OUT[14]_i_2__2 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[30]),
        .I2(crc_from_8[26]),
        .O(\CRC_OUT[14]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \CRC_OUT[14]_i_3__0 
       (.I0(crc_from_8[27]),
        .I1(\CRC_OUT_reg[30]_0 [3]),
        .I2(\CRC_OUT_reg[30]_0 [7]),
        .I3(\CRC_OUT_reg[30]_0 [6]),
        .I4(crc_from_8[6]),
        .O(\CRC_OUT[14]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[15]_i_1__0 
       (.I0(\CRC_OUT[15]_i_2__0_n_0 ),
        .I1(crc_from_8[29]),
        .I2(crc_from_8[31]),
        .I3(\CRC_OUT[15]_i_3__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [15]),
        .O(p_1_in[15]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[15]_i_2__0 
       (.I0(crc_from_8[28]),
        .I1(crc_from_8[27]),
        .O(\CRC_OUT[15]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[15]_i_3__0 
       (.I0(\CRC_OUT_reg[30]_0 [5]),
        .I1(\CRC_OUT_reg[30]_0 [4]),
        .I2(\CRC_OUT_reg[30]_0 [7]),
        .I3(crc_from_8[7]),
        .I4(\CRC_OUT_reg[30]_0 [3]),
        .O(\CRC_OUT[15]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[16]_i_1__0 
       (.I0(\CRC_OUT[16]_i_2__0_n_0 ),
        .I1(crc_from_8[8]),
        .I2(\CRC_OUT[16]_i_3__0_n_0 ),
        .I3(\CRC_OUT[16]_i_4__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [16]),
        .O(p_1_in[16]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[16]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [0]),
        .I1(crc_from_8[24]),
        .O(\CRC_OUT[16]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[16]_i_3__0 
       (.I0(crc_from_8[29]),
        .I1(crc_from_8[28]),
        .O(\CRC_OUT[16]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[16]_i_4__0 
       (.I0(\CRC_OUT_reg[30]_0 [5]),
        .I1(\CRC_OUT_reg[30]_0 [4]),
        .O(\CRC_OUT[16]_i_4__0_n_0 ));
  LUT4 #(
    .INIT(16'h6F60)) 
    \CRC_OUT[17]_i_1__0 
       (.I0(crc_from_8[30]),
        .I1(\CRC_OUT[17]_i_2__0_n_0 ),
        .I2(\CRC_OUT_reg[19]_0 ),
        .I3(\CRC_OUT_reg[31]_0 [17]),
        .O(p_1_in[17]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [6]),
        .I1(\CRC_OUT_reg[30]_0 [5]),
        .I2(crc_from_8[9]),
        .I3(crc_from_8[25]),
        .I4(\CRC_OUT_reg[30]_0 [1]),
        .I5(crc_from_8[29]),
        .O(\CRC_OUT[17]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[18]_i_1__0 
       (.I0(crc_from_8[30]),
        .I1(\CRC_OUT[18]_i_2__1_n_0 ),
        .I2(crc_from_8[10]),
        .I3(\CRC_OUT[18]_i_3__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [18]),
        .O(p_1_in[18]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \CRC_OUT[18]_i_2__1 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(\CRC_OUT_reg[30]_0 [6]),
        .I2(\CRC_OUT_reg[30]_0 [7]),
        .O(\CRC_OUT[18]_i_2__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_3__0 
       (.I0(crc_from_8[26]),
        .I1(crc_from_8[31]),
        .O(\CRC_OUT[18]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[19]_i_1__0 
       (.I0(crc_from_8[27]),
        .I1(crc_from_8[31]),
        .I2(\CRC_OUT[19]_i_2__0_n_0 ),
        .I3(crc_from_8[11]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [19]),
        .O(p_1_in[19]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[19]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [7]),
        .I1(\CRC_OUT_reg[30]_0 [3]),
        .O(\CRC_OUT[19]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[1]_i_1__0 
       (.I0(\CRC_OUT[23]_i_2__0_n_0 ),
        .I1(crc_from_8[30]),
        .I2(crc_from_8[31]),
        .I3(\CRC_OUT[13]_i_3__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [1]),
        .O(p_1_in[1]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[20]_i_1__0 
       (.I0(crc_from_8[12]),
        .I1(crc_from_8[28]),
        .I2(\CRC_OUT_reg[30]_0 [4]),
        .I3(\CRC_OUT_reg[19]_0 ),
        .I4(\CRC_OUT_reg[31]_0 [20]),
        .O(p_1_in[20]));
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[21]_i_1__0 
       (.I0(crc_from_8[13]),
        .I1(crc_from_8[29]),
        .I2(\CRC_OUT_reg[30]_0 [5]),
        .I3(\CRC_OUT_reg[19]_0 ),
        .I4(\CRC_OUT_reg[31]_0 [21]),
        .O(p_1_in[21]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[22]_i_1__0 
       (.I0(crc_from_8[14]),
        .I1(crc_from_8[24]),
        .I2(\CRC_OUT_reg[30]_0 [0]),
        .I3(\CRC_OUT_reg[19]_0 ),
        .I4(\CRC_OUT_reg[31]_0 [22]),
        .O(p_1_in[22]));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[23]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [6]),
        .I1(crc_from_8[30]),
        .I2(crc_from_8[15]),
        .I3(\CRC_OUT[23]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [23]),
        .O(p_1_in[23]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[23]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [1]),
        .I1(crc_from_8[25]),
        .I2(crc_from_8[24]),
        .I3(\CRC_OUT_reg[30]_0 [0]),
        .O(\CRC_OUT[23]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[24]_i_1__0 
       (.I0(\CRC_OUT[24]_i_2__0_n_0 ),
        .I1(crc_from_8[16]),
        .I2(\CRC_OUT[24]_i_3__0_n_0 ),
        .I3(\CRC_OUT[24]_i_4__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [24]),
        .O(p_1_in[24]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [7]),
        .I1(crc_from_8[31]),
        .O(\CRC_OUT[24]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_3__0 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[26]),
        .O(\CRC_OUT[24]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_4__0 
       (.I0(crc_from_8[25]),
        .I1(\CRC_OUT_reg[30]_0 [1]),
        .O(\CRC_OUT[24]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[25]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [3]),
        .I1(\CRC_OUT_reg[30]_0 [2]),
        .I2(\CRC_OUT[25]_i_2__0_n_0 ),
        .I3(crc_from_8[17]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [25]),
        .O(p_1_in[25]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_2__0 
       (.I0(crc_from_8[26]),
        .I1(crc_from_8[27]),
        .O(\CRC_OUT[25]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[26]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [6]),
        .I1(\CRC_OUT_reg[30]_0 [3]),
        .I2(\CRC_OUT_reg[30]_0 [4]),
        .I3(\CRC_OUT[26]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [26]),
        .O(p_1_in[26]));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[26]_i_2__0 
       (.I0(crc_from_8[28]),
        .I1(crc_from_8[27]),
        .I2(crc_from_8[18]),
        .I3(\CRC_OUT_reg[30]_0 [0]),
        .I4(crc_from_8[24]),
        .I5(crc_from_8[30]),
        .O(\CRC_OUT[26]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[27]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [5]),
        .I1(\CRC_OUT_reg[30]_0 [4]),
        .I2(\CRC_OUT_reg[30]_0 [7]),
        .I3(\CRC_OUT[27]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [27]),
        .O(p_1_in[27]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_2__0 
       (.I0(crc_from_8[25]),
        .I1(\CRC_OUT_reg[30]_0 [1]),
        .I2(crc_from_8[19]),
        .I3(crc_from_8[29]),
        .I4(crc_from_8[28]),
        .I5(crc_from_8[31]),
        .O(\CRC_OUT[27]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[28]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[29]),
        .I2(crc_from_8[20]),
        .I3(\CRC_OUT[28]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [28]),
        .O(p_1_in[28]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [5]),
        .I1(\CRC_OUT_reg[30]_0 [6]),
        .I2(crc_from_8[30]),
        .I3(crc_from_8[26]),
        .O(\CRC_OUT[28]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[29]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [7]),
        .I1(\CRC_OUT_reg[30]_0 [6]),
        .I2(crc_from_8[21]),
        .I3(\CRC_OUT[29]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [29]),
        .O(p_1_in[29]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[29]_i_2__0 
       (.I0(crc_from_8[27]),
        .I1(crc_from_8[31]),
        .I2(crc_from_8[30]),
        .I3(\CRC_OUT_reg[30]_0 [3]),
        .O(\CRC_OUT[29]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[2]_i_1__0 
       (.I0(\CRC_OUT[2]_i_2__0_n_0 ),
        .I1(\CRC_OUT_reg[30]_0 [2]),
        .I2(\CRC_OUT[13]_i_3__0_n_0 ),
        .I3(\CRC_OUT[16]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [2]),
        .O(p_1_in[2]));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \CRC_OUT[2]_i_2__0 
       (.I0(crc_from_8[25]),
        .I1(\CRC_OUT_reg[30]_0 [1]),
        .I2(crc_from_8[30]),
        .I3(crc_from_8[31]),
        .I4(crc_from_8[26]),
        .O(\CRC_OUT[2]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[30]_i_1__0 
       (.I0(crc_from_8[31]),
        .I1(\CRC_OUT_reg[30]_0 [7]),
        .I2(\CRC_OUT[30]_i_2__0_n_0 ),
        .I3(crc_from_8[22]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [30]),
        .O(p_1_in[30]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[30]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [4]),
        .I1(crc_from_8[28]),
        .O(\CRC_OUT[30]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \CRC_OUT[31]_i_1 
       (.I0(crc_from_8[23]),
        .I1(crc_from_8[29]),
        .I2(\CRC_OUT_reg[30]_0 [5]),
        .I3(\CRC_OUT_reg[19]_0 ),
        .I4(\CRC_OUT_reg[31]_0 [31]),
        .O(p_1_in[31]));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[3]_i_1__0 
       (.I0(\CRC_OUT[24]_i_3__0_n_0 ),
        .I1(\CRC_OUT[3]_i_2__2_n_0 ),
        .I2(\CRC_OUT[19]_i_2__0_n_0 ),
        .I3(\CRC_OUT[24]_i_4__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [3]),
        .O(p_1_in[3]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \CRC_OUT[3]_i_2__2 
       (.I0(crc_from_8[31]),
        .I1(crc_from_8[27]),
        .O(\CRC_OUT[3]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[4]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [6]),
        .I1(\CRC_OUT_reg[30]_0 [3]),
        .I2(\CRC_OUT_reg[30]_0 [4]),
        .I3(\CRC_OUT[4]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [4]),
        .O(p_1_in[4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_2__0 
       (.I0(\CRC_OUT[16]_i_2__0_n_0 ),
        .I1(\CRC_OUT_reg[30]_0 [2]),
        .I2(crc_from_8[28]),
        .I3(crc_from_8[27]),
        .I4(crc_from_8[26]),
        .I5(crc_from_8[30]),
        .O(\CRC_OUT[4]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[5]_i_1__0 
       (.I0(\CRC_OUT[23]_i_2__0_n_0 ),
        .I1(crc_from_8[28]),
        .I2(crc_from_8[27]),
        .I3(\CRC_OUT[5]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [5]),
        .O(p_1_in[5]));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[5]_i_2__0 
       (.I0(crc_from_8[29]),
        .I1(crc_from_8[31]),
        .I2(crc_from_8[30]),
        .I3(\CRC_OUT[5]_i_3__1_n_0 ),
        .I4(\CRC_OUT_reg[30]_0 [7]),
        .I5(\CRC_OUT_reg[30]_0 [5]),
        .O(\CRC_OUT[5]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \CRC_OUT[5]_i_3__1 
       (.I0(\CRC_OUT_reg[30]_0 [4]),
        .I1(\CRC_OUT_reg[30]_0 [3]),
        .I2(\CRC_OUT_reg[30]_0 [6]),
        .O(\CRC_OUT[5]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h9669FFFF96690000)) 
    \CRC_OUT[6]_i_1__0 
       (.I0(\CRC_OUT[6]_i_2__0_n_0 ),
        .I1(\CRC_OUT_reg[30]_0 [5]),
        .I2(\CRC_OUT[13]_i_3__0_n_0 ),
        .I3(\CRC_OUT[24]_i_4__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [6]),
        .O(p_1_in[6]));
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \CRC_OUT[6]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[30]),
        .I2(\CRC_OUT_reg[30]_0 [4]),
        .I3(crc_from_8[26]),
        .I4(crc_from_8[31]),
        .I5(\CRC_OUT[16]_i_3__0_n_0 ),
        .O(\CRC_OUT[6]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[7]_i_1__0 
       (.I0(\CRC_OUT[25]_i_2__0_n_0 ),
        .I1(crc_from_8[29]),
        .I2(crc_from_8[31]),
        .I3(\CRC_OUT[7]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [7]),
        .O(p_1_in[7]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[7]_i_2__0 
       (.I0(\CRC_OUT_reg[30]_0 [0]),
        .I1(crc_from_8[24]),
        .I2(\CRC_OUT_reg[30]_0 [2]),
        .I3(\CRC_OUT_reg[30]_0 [7]),
        .I4(\CRC_OUT_reg[30]_0 [3]),
        .I5(\CRC_OUT_reg[30]_0 [5]),
        .O(\CRC_OUT[7]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[8]_i_1__0 
       (.I0(crc_from_8[0]),
        .I1(\CRC_OUT[11]_i_2__0_n_0 ),
        .I2(\CRC_OUT_reg[30]_0 [3]),
        .I3(\CRC_OUT_reg[30]_0 [4]),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [8]),
        .O(p_1_in[8]));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \CRC_OUT[9]_i_1__0 
       (.I0(\CRC_OUT_reg[30]_0 [2]),
        .I1(crc_from_8[26]),
        .I2(\CRC_OUT[16]_i_3__0_n_0 ),
        .I3(\CRC_OUT[9]_i_2__0_n_0 ),
        .I4(\CRC_OUT_reg[19]_0 ),
        .I5(\CRC_OUT_reg[31]_0 [9]),
        .O(p_1_in[9]));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[9]_i_2__0 
       (.I0(crc_from_8[1]),
        .I1(crc_from_8[25]),
        .I2(\CRC_OUT_reg[30]_0 [1]),
        .I3(\CRC_OUT_reg[30]_0 [5]),
        .I4(\CRC_OUT_reg[30]_0 [4]),
        .O(\CRC_OUT[9]_i_2__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[0]),
        .Q(crc_from_8[0]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[10]),
        .Q(crc_from_8[10]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[11]),
        .Q(crc_from_8[11]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[12]),
        .Q(crc_from_8[12]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[13]),
        .Q(crc_from_8[13]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[14]),
        .Q(crc_from_8[14]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[15]),
        .Q(crc_from_8[15]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[16]),
        .Q(crc_from_8[16]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[17]),
        .Q(crc_from_8[17]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[18]),
        .Q(crc_from_8[18]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[19]),
        .Q(crc_from_8[19]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[1]),
        .Q(crc_from_8[1]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[20]),
        .Q(crc_from_8[20]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[21]),
        .Q(crc_from_8[21]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[22]),
        .Q(crc_from_8[22]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[23]),
        .Q(crc_from_8[23]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[24]),
        .Q(crc_from_8[24]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[25]),
        .Q(crc_from_8[25]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[26]),
        .Q(crc_from_8[26]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[27]),
        .Q(crc_from_8[27]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[28]),
        .Q(crc_from_8[28]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[29]),
        .Q(crc_from_8[29]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[2]),
        .Q(crc_from_8[2]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[30]),
        .Q(crc_from_8[30]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[31]),
        .Q(crc_from_8[31]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[3]),
        .Q(crc_from_8[3]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[4]),
        .Q(crc_from_8[4]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[5]),
        .Q(crc_from_8[5]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[6]),
        .Q(crc_from_8[6]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[7]),
        .Q(crc_from_8[7]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[8]),
        .Q(crc_from_8[8]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_OUT_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_1_in[9]),
        .Q(crc_from_8[9]));
  LUT5 #(
    .INIT(32'h00000002)) 
    good_frame_get_i_2
       (.I0(good_frame_get_i_3_n_0),
        .I1(D),
        .I2(small_error),
        .I3(large_error),
        .I4(Q),
        .O(small_error_reg));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    good_frame_get_i_3
       (.I0(\rxStatRegPlus[1]_i_2_n_0 ),
        .I1(\rxStatRegPlus[1]_i_5_n_0 ),
        .I2(\rxStatRegPlus[1]_i_4_n_0 ),
        .I3(do_crc_check),
        .I4(wait_crc_check),
        .I5(\rxStatRegPlus[1]_i_3_n_0 ),
        .O(good_frame_get_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFD000000000000)) 
    \rxStatRegPlus[1]_i_1 
       (.I0(\rxStatRegPlus[1]_i_2_n_0 ),
        .I1(\rxStatRegPlus[1]_i_3_n_0 ),
        .I2(\rxStatRegPlus[1]_i_4_n_0 ),
        .I3(\rxStatRegPlus[1]_i_5_n_0 ),
        .I4(wait_crc_check),
        .I5(do_crc_check),
        .O(D));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \rxStatRegPlus[1]_i_10 
       (.I0(crc_from_8[1]),
        .I1(crc_from_8[16]),
        .I2(crc_from_8[21]),
        .I3(crc_from_8[20]),
        .O(\rxStatRegPlus[1]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \rxStatRegPlus[1]_i_2 
       (.I0(\rxStatRegPlus[1]_i_6_n_0 ),
        .I1(\rxStatRegPlus[1]_i_7_n_0 ),
        .I2(\rxStatRegPlus[1]_i_8_n_0 ),
        .I3(\rxStatRegPlus[1]_i_9_n_0 ),
        .I4(\rxStatRegPlus[1]_i_10_n_0 ),
        .O(\rxStatRegPlus[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF7)) 
    \rxStatRegPlus[1]_i_3 
       (.I0(crc_from_8[11]),
        .I1(crc_from_8[10]),
        .I2(crc_from_8[7]),
        .I3(crc_from_8[9]),
        .I4(crc_from_8[13]),
        .O(\rxStatRegPlus[1]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \rxStatRegPlus[1]_i_4 
       (.I0(crc_from_8[29]),
        .I1(crc_from_8[27]),
        .I2(crc_from_8[28]),
        .O(\rxStatRegPlus[1]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rxStatRegPlus[1]_i_5 
       (.I0(crc_from_8[5]),
        .I1(crc_from_8[4]),
        .I2(crc_from_8[31]),
        .I3(crc_from_8[30]),
        .O(\rxStatRegPlus[1]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rxStatRegPlus[1]_i_6 
       (.I0(crc_from_8[18]),
        .I1(crc_from_8[26]),
        .I2(crc_from_8[12]),
        .I3(crc_from_8[25]),
        .O(\rxStatRegPlus[1]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \rxStatRegPlus[1]_i_7 
       (.I0(crc_from_8[17]),
        .I1(crc_from_8[8]),
        .I2(crc_from_8[6]),
        .I3(crc_from_8[22]),
        .O(\rxStatRegPlus[1]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \rxStatRegPlus[1]_i_8 
       (.I0(crc_from_8[0]),
        .I1(crc_from_8[19]),
        .I2(crc_from_8[15]),
        .I3(crc_from_8[14]),
        .O(\rxStatRegPlus[1]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hFFDF)) 
    \rxStatRegPlus[1]_i_9 
       (.I0(crc_from_8[3]),
        .I1(crc_from_8[23]),
        .I2(crc_from_8[24]),
        .I3(crc_from_8[2]),
        .O(\rxStatRegPlus[1]_i_9_n_0 ));
endmodule

(* ORIG_REF_NAME = "Calculator" *) 
module switch_elements_Calculator
   (D,
    \A0_reg[11]_0 ,
    Q,
    \B1_reg[11]_0 ,
    \t3z3_reg[18] ,
    doii1,
    \shii_reg[0]_0 ,
    \d1_4_reg[15] ,
    \d2_4_reg[15] ,
    \d3_4_reg[15] ,
    \a0d_reg[11] ,
    O,
    \z1d1_reg[15] ,
    \z1d1_reg[15]_0 ,
    \z1d1_reg[15]_1 ,
    \z1d1_reg[15]_2 ,
    \z2d1_reg[15] ,
    \z2d1_reg[15]_0 ,
    \z2d1_reg[15]_1 ,
    \z2d1_reg[15]_2 ,
    \z3d1_reg[15] ,
    \z3d1_reg[15]_0 ,
    \z3d1_reg[15]_1 ,
    \z3d1_reg[15]_2 ,
    FREQ,
    clk_i,
    rst_i,
    out);
  output [11:0]D;
  output [11:0]\A0_reg[11]_0 ;
  output [0:0]Q;
  output [11:0]\B1_reg[11]_0 ;
  output [1:0]\t3z3_reg[18] ;
  output doii1;
  output \shii_reg[0]_0 ;
  output [15:0]\d1_4_reg[15] ;
  output [15:0]\d2_4_reg[15] ;
  output [15:0]\d3_4_reg[15] ;
  input [2:0]\a0d_reg[11] ;
  input [1:0]O;
  input [15:0]\z1d1_reg[15] ;
  input [15:0]\z1d1_reg[15]_0 ;
  input [15:0]\z1d1_reg[15]_1 ;
  input [15:0]\z1d1_reg[15]_2 ;
  input [15:0]\z2d1_reg[15] ;
  input [15:0]\z2d1_reg[15]_0 ;
  input [15:0]\z2d1_reg[15]_1 ;
  input [15:0]\z2d1_reg[15]_2 ;
  input [15:0]\z3d1_reg[15] ;
  input [15:0]\z3d1_reg[15]_0 ;
  input [15:0]\z3d1_reg[15]_1 ;
  input [15:0]\z3d1_reg[15]_2 ;
  input [11:0]FREQ;
  input clk_i;
  input rst_i;
  input out;

  wire [11:0]A0;
  wire [11:0]\A0_reg[11]_0 ;
  wire [11:0]A1;
  wire [11:0]B1;
  wire [11:0]\B1_reg[11]_0 ;
  wire [11:0]D;
  wire [11:0]FREQ;
  wire [1:0]O;
  wire [0:0]Q;
  wire \_inferred__4/i__carry__0_n_5 ;
  wire \_inferred__4/i__carry__0_n_6 ;
  wire \_inferred__4/i__carry__0_n_7 ;
  wire \_inferred__4/i__carry_n_0 ;
  wire \_inferred__4/i__carry_n_1 ;
  wire \_inferred__4/i__carry_n_2 ;
  wire \_inferred__4/i__carry_n_3 ;
  wire \_inferred__4/i__carry_n_4 ;
  wire \_inferred__4/i__carry_n_5 ;
  wire \_inferred__4/i__carry_n_6 ;
  wire \_inferred__4/i__carry_n_7 ;
  wire [11:0]a;
  wire [2:0]\a0d_reg[11] ;
  wire a11;
  wire a_0;
  wire b11;
  wire \b1d[11]_i_3_n_0 ;
  wire clk_i;
  wire [15:0]\d1_4_reg[15] ;
  wire [15:0]\d2_4_reg[15] ;
  wire [15:0]\d3_4_reg[15] ;
  wire doii1;
  wire ea0;
  wire ea1;
  wire eb1;
  wire esh;
  wire [11:0]fi;
  wire g0_b0__0__0_n_0;
  wire g0_b0__0_n_0;
  wire g0_b0__10_n_0;
  wire g0_b0__1_n_0;
  wire g0_b0__2_n_0;
  wire g0_b0__3_n_0;
  wire g0_b0__4_n_0;
  wire g0_b0__5_n_0;
  wire g0_b0__6_n_0;
  wire g0_b0__7_n_0;
  wire g0_b0__8_n_0;
  wire g0_b0__9_n_0;
  wire g0_b0_n_0;
  wire i__carry__0_i_4_n_0;
  wire i__carry__0_i_5_n_0;
  wire i__carry__0_i_6_n_0;
  wire i__carry__0_i_7_n_0;
  wire i__carry_i_10__2_n_0;
  wire i__carry_i_11__4_n_0;
  wire i__carry_i_12__0_n_0;
  wire i__carry_i_13_n_0;
  wire i__carry_i_14_n_0;
  wire i__carry_i_15_n_0;
  wire i__carry_i_16_n_0;
  wire i__carry_i_17_n_0;
  wire i__carry_i_18_n_0;
  wire i__carry_i_19_n_0;
  wire i__carry_i_1__2_n_0;
  wire i__carry_i_20_n_0;
  wire i__carry_i_21_n_0;
  wire i__carry_i_22_n_0;
  wire i__carry_i_23_n_0;
  wire i__carry_i_24_n_0;
  wire i__carry_i_25_n_0;
  wire i__carry_i_26_n_0;
  wire i__carry_i_27_n_0;
  wire i__carry_i_28_n_0;
  wire i__carry_i_29_n_0;
  wire i__carry_i_30_n_0;
  wire i__carry_i_31_n_0;
  wire i__carry_i_32_n_0;
  wire i__carry_i_33_n_0;
  wire i__carry_i_34_n_0;
  wire i__carry_i_35_n_0;
  wire out;
  wire [10:1]p_1_in__1;
  wire p_2_in;
  wire [4:0]plusOp__0;
  wire [11:0]q;
  wire rst_i;
  wire [2:1]sel0;
  wire [3:1]sh;
  wire [3:1]shi;
  wire \shii[0]_i_1_n_0 ;
  wire \shii_reg[0]_0 ;
  wire [11:0]sr;
  wire \sr[0]_i_1_n_0 ;
  wire \sr[10]_i_1_n_0 ;
  wire \sr[10]_i_2_n_0 ;
  wire \sr[10]_i_3_n_0 ;
  wire \sr[11]_i_1_n_0 ;
  wire \sr[1]_i_1_n_0 ;
  wire \sr[2]_i_1_n_0 ;
  wire \sr[3]_i_1_n_0 ;
  wire \sr[4]_i_1_n_0 ;
  wire \sr[5]_i_1_n_0 ;
  wire \sr[6]_i_1_n_0 ;
  wire \sr[7]_i_1_n_0 ;
  wire \sr[8]_i_1_n_0 ;
  wire \sr[9]_i_1_n_0 ;
  wire \st[3]_i_1_n_0 ;
  wire \st[4]_i_1_n_0 ;
  wire [4:0]st_reg;
  wire [1:0]\t3z3_reg[18] ;
  wire [15:0]\z1d1_reg[15] ;
  wire [15:0]\z1d1_reg[15]_0 ;
  wire [15:0]\z1d1_reg[15]_1 ;
  wire [15:0]\z1d1_reg[15]_2 ;
  wire [15:0]\z2d1_reg[15] ;
  wire [15:0]\z2d1_reg[15]_0 ;
  wire [15:0]\z2d1_reg[15]_1 ;
  wire [15:0]\z2d1_reg[15]_2 ;
  wire [15:0]\z3d1_reg[15] ;
  wire [15:0]\z3d1_reg[15]_0 ;
  wire [15:0]\z3d1_reg[15]_1 ;
  wire [15:0]\z3d1_reg[15]_2 ;
  wire [7:3]\NLW__inferred__4/i__carry__0_CO_UNCONNECTED ;
  wire [7:4]\NLW__inferred__4/i__carry__0_O_UNCONNECTED ;

  LUT5 #(
    .INIT(32'h00001000)) 
    \A0[11]_i_1 
       (.I0(st_reg[2]),
        .I1(st_reg[3]),
        .I2(st_reg[4]),
        .I3(st_reg[0]),
        .I4(st_reg[1]),
        .O(ea0));
  FDCE #(
    .INIT(1'b0)) 
    \A0_reg[0] 
       (.C(clk_i),
        .CE(ea0),
        .CLR(rst_i),
        .D(q[0]),
        .Q(A0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \A0_reg[10] 
       (.C(clk_i),
        .CE(ea0),
        .CLR(rst_i),
        .D(q[10]),
        .Q(A0[10]));
  FDCE #(
    .INIT(1'b0)) 
    \A0_reg[11] 
       (.C(clk_i),
        .CE(ea0),
        .CLR(rst_i),
        .D(q[11]),
        .Q(A0[11]));
  FDCE #(
    .INIT(1'b0)) 
    \A0_reg[1] 
       (.C(clk_i),
        .CE(ea0),
        .CLR(rst_i),
        .D(q[1]),
        .Q(A0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \A0_reg[2] 
       (.C(clk_i),
        .CE(ea0),
        .CLR(rst_i),
        .D(q[2]),
        .Q(A0[2]));
  FDPE #(
    .INIT(1'b1)) 
    \A0_reg[3] 
       (.C(clk_i),
        .CE(ea0),
        .D(q[3]),
        .PRE(rst_i),
        .Q(A0[3]));
  FDPE #(
    .INIT(1'b1)) 
    \A0_reg[4] 
       (.C(clk_i),
        .CE(ea0),
        .D(q[4]),
        .PRE(rst_i),
        .Q(A0[4]));
  FDPE #(
    .INIT(1'b1)) 
    \A0_reg[5] 
       (.C(clk_i),
        .CE(ea0),
        .D(q[5]),
        .PRE(rst_i),
        .Q(A0[5]));
  FDPE #(
    .INIT(1'b1)) 
    \A0_reg[6] 
       (.C(clk_i),
        .CE(ea0),
        .D(q[6]),
        .PRE(rst_i),
        .Q(A0[6]));
  FDPE #(
    .INIT(1'b1)) 
    \A0_reg[7] 
       (.C(clk_i),
        .CE(ea0),
        .D(q[7]),
        .PRE(rst_i),
        .Q(A0[7]));
  FDPE #(
    .INIT(1'b1)) 
    \A0_reg[8] 
       (.C(clk_i),
        .CE(ea0),
        .D(q[8]),
        .PRE(rst_i),
        .Q(A0[8]));
  FDCE #(
    .INIT(1'b0)) 
    \A0_reg[9] 
       (.C(clk_i),
        .CE(ea0),
        .CLR(rst_i),
        .D(q[9]),
        .Q(A0[9]));
  LUT5 #(
    .INIT(32'h00100000)) 
    \A1[11]_i_1 
       (.I0(st_reg[4]),
        .I1(st_reg[2]),
        .I2(st_reg[3]),
        .I3(st_reg[1]),
        .I4(st_reg[0]),
        .O(ea1));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[0] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[0]),
        .PRE(rst_i),
        .Q(A1[0]));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[10] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[10]),
        .PRE(rst_i),
        .Q(A1[10]));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[11] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[11]),
        .PRE(rst_i),
        .Q(A1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \A1_reg[1] 
       (.C(clk_i),
        .CE(ea1),
        .CLR(rst_i),
        .D(q[1]),
        .Q(A1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \A1_reg[2] 
       (.C(clk_i),
        .CE(ea1),
        .CLR(rst_i),
        .D(q[2]),
        .Q(A1[2]));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[3] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[3]),
        .PRE(rst_i),
        .Q(A1[3]));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[4] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[4]),
        .PRE(rst_i),
        .Q(A1[4]));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[5] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[5]),
        .PRE(rst_i),
        .Q(A1[5]));
  FDPE #(
    .INIT(1'b1)) 
    \A1_reg[6] 
       (.C(clk_i),
        .CE(ea1),
        .D(q[6]),
        .PRE(rst_i),
        .Q(A1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \A1_reg[7] 
       (.C(clk_i),
        .CE(ea1),
        .CLR(rst_i),
        .D(q[7]),
        .Q(A1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \A1_reg[8] 
       (.C(clk_i),
        .CE(ea1),
        .CLR(rst_i),
        .D(q[8]),
        .Q(A1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \A1_reg[9] 
       (.C(clk_i),
        .CE(ea1),
        .CLR(rst_i),
        .D(q[9]),
        .Q(A1[9]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \B1[11]_i_1 
       (.I0(st_reg[4]),
        .I1(st_reg[3]),
        .I2(st_reg[0]),
        .I3(st_reg[2]),
        .I4(st_reg[1]),
        .O(eb1));
  FDPE #(
    .INIT(1'b1)) 
    \B1_reg[0] 
       (.C(clk_i),
        .CE(eb1),
        .D(q[0]),
        .PRE(rst_i),
        .Q(B1[0]));
  FDPE #(
    .INIT(1'b1)) 
    \B1_reg[10] 
       (.C(clk_i),
        .CE(eb1),
        .D(q[10]),
        .PRE(rst_i),
        .Q(B1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[11] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[11]),
        .Q(B1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[1] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[1]),
        .Q(B1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[2] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[2]),
        .Q(B1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[3] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[3]),
        .Q(B1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[4] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[4]),
        .Q(B1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[5] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[5]),
        .Q(B1[5]));
  FDPE #(
    .INIT(1'b1)) 
    \B1_reg[6] 
       (.C(clk_i),
        .CE(eb1),
        .D(q[6]),
        .PRE(rst_i),
        .Q(B1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[7] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[7]),
        .Q(B1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[8] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[8]),
        .Q(B1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \B1_reg[9] 
       (.C(clk_i),
        .CE(eb1),
        .CLR(rst_i),
        .D(q[9]),
        .Q(B1[9]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[0].U_SRL_i_1__2 
       (.I0(\z1d1_reg[15] [0]),
        .I1(\z1d1_reg[15]_0 [0]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [0]),
        .I5(\z1d1_reg[15]_2 [0]),
        .O(\d1_4_reg[15] [0]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[0].U_SRL_i_1__3 
       (.I0(\z2d1_reg[15] [0]),
        .I1(\z2d1_reg[15]_0 [0]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [0]),
        .I5(\z2d1_reg[15]_2 [0]),
        .O(\d2_4_reg[15] [0]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[0].U_SRL_i_1__4 
       (.I0(\z3d1_reg[15] [0]),
        .I1(\z3d1_reg[15]_0 [0]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [0]),
        .I5(\z3d1_reg[15]_2 [0]),
        .O(\d3_4_reg[15] [0]));
  LUT6 #(
    .INIT(64'h3CCC2CC83CCC2888)) 
    \D16.DEL0[0].U_SRL_i_2 
       (.I0(Q),
        .I1(\a0d_reg[11] [2]),
        .I2(\a0d_reg[11] [0]),
        .I3(\a0d_reg[11] [1]),
        .I4(sh[1]),
        .I5(sh[2]),
        .O(doii1));
  LUT3 #(
    .INIT(8'hF4)) 
    \D16.DEL0[0].U_SRL_i_2__0 
       (.I0(\a0d_reg[11] [2]),
        .I1(Q),
        .I2(\a0d_reg[11] [1]),
        .O(sel0[1]));
  LUT3 #(
    .INIT(8'hF4)) 
    \D16.DEL0[0].U_SRL_i_3 
       (.I0(\a0d_reg[11] [1]),
        .I1(Q),
        .I2(\a0d_reg[11] [2]),
        .O(sel0[2]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[10].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [10]),
        .I1(\z1d1_reg[15]_0 [10]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [10]),
        .I5(\z1d1_reg[15]_2 [10]),
        .O(\d1_4_reg[15] [10]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[10].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [10]),
        .I1(\z2d1_reg[15]_0 [10]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [10]),
        .I5(\z2d1_reg[15]_2 [10]),
        .O(\d2_4_reg[15] [10]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[10].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [10]),
        .I1(\z3d1_reg[15]_0 [10]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [10]),
        .I5(\z3d1_reg[15]_2 [10]),
        .O(\d3_4_reg[15] [10]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[11].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [11]),
        .I1(\z1d1_reg[15]_0 [11]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [11]),
        .I5(\z1d1_reg[15]_2 [11]),
        .O(\d1_4_reg[15] [11]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[11].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [11]),
        .I1(\z2d1_reg[15]_0 [11]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [11]),
        .I5(\z2d1_reg[15]_2 [11]),
        .O(\d2_4_reg[15] [11]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[11].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [11]),
        .I1(\z3d1_reg[15]_0 [11]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [11]),
        .I5(\z3d1_reg[15]_2 [11]),
        .O(\d3_4_reg[15] [11]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[12].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [12]),
        .I1(\z1d1_reg[15]_0 [12]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [12]),
        .I5(\z1d1_reg[15]_2 [12]),
        .O(\d1_4_reg[15] [12]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[12].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [12]),
        .I1(\z2d1_reg[15]_0 [12]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [12]),
        .I5(\z2d1_reg[15]_2 [12]),
        .O(\d2_4_reg[15] [12]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[12].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [12]),
        .I1(\z3d1_reg[15]_0 [12]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [12]),
        .I5(\z3d1_reg[15]_2 [12]),
        .O(\d3_4_reg[15] [12]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[13].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [13]),
        .I1(\z1d1_reg[15]_0 [13]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [13]),
        .I5(\z1d1_reg[15]_2 [13]),
        .O(\d1_4_reg[15] [13]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[13].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [13]),
        .I1(\z2d1_reg[15]_0 [13]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [13]),
        .I5(\z2d1_reg[15]_2 [13]),
        .O(\d2_4_reg[15] [13]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[13].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [13]),
        .I1(\z3d1_reg[15]_0 [13]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [13]),
        .I5(\z3d1_reg[15]_2 [13]),
        .O(\d3_4_reg[15] [13]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[14].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [14]),
        .I1(\z1d1_reg[15]_0 [14]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [14]),
        .I5(\z1d1_reg[15]_2 [14]),
        .O(\d1_4_reg[15] [14]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[14].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [14]),
        .I1(\z2d1_reg[15]_0 [14]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [14]),
        .I5(\z2d1_reg[15]_2 [14]),
        .O(\d2_4_reg[15] [14]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[14].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [14]),
        .I1(\z3d1_reg[15]_0 [14]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [14]),
        .I5(\z3d1_reg[15]_2 [14]),
        .O(\d3_4_reg[15] [14]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[15].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [15]),
        .I1(\z1d1_reg[15]_0 [15]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [15]),
        .I5(\z1d1_reg[15]_2 [15]),
        .O(\d1_4_reg[15] [15]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[15].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [15]),
        .I1(\z2d1_reg[15]_0 [15]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [15]),
        .I5(\z2d1_reg[15]_2 [15]),
        .O(\d2_4_reg[15] [15]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[15].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [15]),
        .I1(\z3d1_reg[15]_0 [15]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [15]),
        .I5(\z3d1_reg[15]_2 [15]),
        .O(\d3_4_reg[15] [15]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[1].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [1]),
        .I1(\z1d1_reg[15]_0 [1]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [1]),
        .I5(\z1d1_reg[15]_2 [1]),
        .O(\d1_4_reg[15] [1]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[1].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [1]),
        .I1(\z2d1_reg[15]_0 [1]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [1]),
        .I5(\z2d1_reg[15]_2 [1]),
        .O(\d2_4_reg[15] [1]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[1].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [1]),
        .I1(\z3d1_reg[15]_0 [1]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [1]),
        .I5(\z3d1_reg[15]_2 [1]),
        .O(\d3_4_reg[15] [1]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[2].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [2]),
        .I1(\z1d1_reg[15]_0 [2]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [2]),
        .I5(\z1d1_reg[15]_2 [2]),
        .O(\d1_4_reg[15] [2]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[2].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [2]),
        .I1(\z2d1_reg[15]_0 [2]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [2]),
        .I5(\z2d1_reg[15]_2 [2]),
        .O(\d2_4_reg[15] [2]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[2].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [2]),
        .I1(\z3d1_reg[15]_0 [2]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [2]),
        .I5(\z3d1_reg[15]_2 [2]),
        .O(\d3_4_reg[15] [2]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[3].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [3]),
        .I1(\z1d1_reg[15]_0 [3]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [3]),
        .I5(\z1d1_reg[15]_2 [3]),
        .O(\d1_4_reg[15] [3]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[3].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [3]),
        .I1(\z2d1_reg[15]_0 [3]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [3]),
        .I5(\z2d1_reg[15]_2 [3]),
        .O(\d2_4_reg[15] [3]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[3].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [3]),
        .I1(\z3d1_reg[15]_0 [3]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [3]),
        .I5(\z3d1_reg[15]_2 [3]),
        .O(\d3_4_reg[15] [3]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[4].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [4]),
        .I1(\z1d1_reg[15]_0 [4]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [4]),
        .I5(\z1d1_reg[15]_2 [4]),
        .O(\d1_4_reg[15] [4]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[4].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [4]),
        .I1(\z2d1_reg[15]_0 [4]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [4]),
        .I5(\z2d1_reg[15]_2 [4]),
        .O(\d2_4_reg[15] [4]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[4].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [4]),
        .I1(\z3d1_reg[15]_0 [4]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [4]),
        .I5(\z3d1_reg[15]_2 [4]),
        .O(\d3_4_reg[15] [4]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[5].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [5]),
        .I1(\z1d1_reg[15]_0 [5]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [5]),
        .I5(\z1d1_reg[15]_2 [5]),
        .O(\d1_4_reg[15] [5]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[5].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [5]),
        .I1(\z2d1_reg[15]_0 [5]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [5]),
        .I5(\z2d1_reg[15]_2 [5]),
        .O(\d2_4_reg[15] [5]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[5].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [5]),
        .I1(\z3d1_reg[15]_0 [5]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [5]),
        .I5(\z3d1_reg[15]_2 [5]),
        .O(\d3_4_reg[15] [5]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[6].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [6]),
        .I1(\z1d1_reg[15]_0 [6]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [6]),
        .I5(\z1d1_reg[15]_2 [6]),
        .O(\d1_4_reg[15] [6]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[6].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [6]),
        .I1(\z2d1_reg[15]_0 [6]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [6]),
        .I5(\z2d1_reg[15]_2 [6]),
        .O(\d2_4_reg[15] [6]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[6].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [6]),
        .I1(\z3d1_reg[15]_0 [6]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [6]),
        .I5(\z3d1_reg[15]_2 [6]),
        .O(\d3_4_reg[15] [6]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[7].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [7]),
        .I1(\z1d1_reg[15]_0 [7]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [7]),
        .I5(\z1d1_reg[15]_2 [7]),
        .O(\d1_4_reg[15] [7]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[7].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [7]),
        .I1(\z2d1_reg[15]_0 [7]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [7]),
        .I5(\z2d1_reg[15]_2 [7]),
        .O(\d2_4_reg[15] [7]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[7].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [7]),
        .I1(\z3d1_reg[15]_0 [7]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [7]),
        .I5(\z3d1_reg[15]_2 [7]),
        .O(\d3_4_reg[15] [7]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[8].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [8]),
        .I1(\z1d1_reg[15]_0 [8]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [8]),
        .I5(\z1d1_reg[15]_2 [8]),
        .O(\d1_4_reg[15] [8]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[8].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [8]),
        .I1(\z2d1_reg[15]_0 [8]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [8]),
        .I5(\z2d1_reg[15]_2 [8]),
        .O(\d2_4_reg[15] [8]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[8].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [8]),
        .I1(\z3d1_reg[15]_0 [8]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [8]),
        .I5(\z3d1_reg[15]_2 [8]),
        .O(\d3_4_reg[15] [8]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[9].U_SRL_i_1__0 
       (.I0(\z1d1_reg[15] [9]),
        .I1(\z1d1_reg[15]_0 [9]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z1d1_reg[15]_1 [9]),
        .I5(\z1d1_reg[15]_2 [9]),
        .O(\d1_4_reg[15] [9]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[9].U_SRL_i_1__1 
       (.I0(\z2d1_reg[15] [9]),
        .I1(\z2d1_reg[15]_0 [9]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z2d1_reg[15]_1 [9]),
        .I5(\z2d1_reg[15]_2 [9]),
        .O(\d2_4_reg[15] [9]));
  LUT6 #(
    .INIT(64'hCFAFCFA0C0AFC0A0)) 
    \D16.DEL0[9].U_SRL_i_1__2 
       (.I0(\z3d1_reg[15] [9]),
        .I1(\z3d1_reg[15]_0 [9]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\z3d1_reg[15]_1 [9]),
        .I5(\z3d1_reg[15]_2 [9]),
        .O(\d3_4_reg[15] [9]));
  LUT4 #(
    .INIT(16'h0440)) 
    \D32.DEL1[0].U_SRL0_i_3 
       (.I0(Q),
        .I1(\a0d_reg[11] [2]),
        .I2(\a0d_reg[11] [0]),
        .I3(\a0d_reg[11] [1]),
        .O(\shii_reg[0]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \DO[14]_i_1 
       (.I0(O[0]),
        .I1(doii1),
        .O(\t3z3_reg[18] [0]));
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \DO[15]_i_2 
       (.I0(O[1]),
        .I1(doii1),
        .O(\t3z3_reg[18] [1]));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \_inferred__4/i__carry 
       (.CI(i__carry_i_1__2_n_0),
        .CI_TOP(1'b0),
        .CO({\_inferred__4/i__carry_n_0 ,\_inferred__4/i__carry_n_1 ,\_inferred__4/i__carry_n_2 ,\_inferred__4/i__carry_n_3 ,\_inferred__4/i__carry_n_4 ,\_inferred__4/i__carry_n_5 ,\_inferred__4/i__carry_n_6 ,\_inferred__4/i__carry_n_7 }),
        .DI({p_1_in__1[7:1],p_2_in}),
        .O(q[7:0]),
        .S({i__carry_i_10__2_n_0,i__carry_i_11__4_n_0,i__carry_i_12__0_n_0,i__carry_i_13_n_0,i__carry_i_14_n_0,i__carry_i_15_n_0,i__carry_i_16_n_0,i__carry_i_17_n_0}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \_inferred__4/i__carry__0 
       (.CI(\_inferred__4/i__carry_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW__inferred__4/i__carry__0_CO_UNCONNECTED [7:3],\_inferred__4/i__carry__0_n_5 ,\_inferred__4/i__carry__0_n_6 ,\_inferred__4/i__carry__0_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,p_1_in__1[10:8]}),
        .O({\NLW__inferred__4/i__carry__0_O_UNCONNECTED [7:4],q[11:8]}),
        .S({1'b0,1'b0,1'b0,1'b0,i__carry__0_i_4_n_0,i__carry__0_i_5_n_0,i__carry__0_i_6_n_0,i__carry__0_i_7_n_0}));
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a0d[0]_i_1 
       (.I0(a11),
        .I1(A0[0]),
        .O(\A0_reg[11]_0 [0]));
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a0d[10]_i_1 
       (.I0(a11),
        .I1(A0[10]),
        .O(\A0_reg[11]_0 [10]));
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a0d[11]_i_1 
       (.I0(a11),
        .I1(A0[11]),
        .O(\A0_reg[11]_0 [11]));
  LUT6 #(
    .INIT(64'hFCFCF0F0FAFAFFF0)) 
    \a0d[11]_i_2 
       (.I0(sh[3]),
        .I1(sh[1]),
        .I2(Q),
        .I3(sh[2]),
        .I4(\a0d_reg[11] [1]),
        .I5(\a0d_reg[11] [2]),
        .O(a11));
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a0d[1]_i_1 
       (.I0(a11),
        .I1(A0[1]),
        .O(\A0_reg[11]_0 [1]));
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a0d[2]_i_1 
       (.I0(a11),
        .I1(A0[2]),
        .O(\A0_reg[11]_0 [2]));
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a0d[3]_i_1 
       (.I0(A0[3]),
        .I1(a11),
        .O(\A0_reg[11]_0 [3]));
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a0d[4]_i_1 
       (.I0(A0[4]),
        .I1(a11),
        .O(\A0_reg[11]_0 [4]));
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a0d[5]_i_1 
       (.I0(A0[5]),
        .I1(a11),
        .O(\A0_reg[11]_0 [5]));
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a0d[6]_i_1 
       (.I0(A0[6]),
        .I1(a11),
        .O(\A0_reg[11]_0 [6]));
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a0d[7]_i_1 
       (.I0(A0[7]),
        .I1(a11),
        .O(\A0_reg[11]_0 [7]));
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a0d[8]_i_1 
       (.I0(A0[8]),
        .I1(a11),
        .O(\A0_reg[11]_0 [8]));
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a0d[9]_i_1 
       (.I0(a11),
        .I1(A0[9]),
        .O(\A0_reg[11]_0 [9]));
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[0]_i_1 
       (.I0(A1[0]),
        .I1(a11),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[10]_i_1 
       (.I0(A1[10]),
        .I1(a11),
        .O(D[10]));
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[11]_i_1 
       (.I0(A1[11]),
        .I1(a11),
        .O(D[11]));
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a1d[1]_i_1 
       (.I0(a11),
        .I1(A1[1]),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a1d[2]_i_1 
       (.I0(a11),
        .I1(A1[2]),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[3]_i_1 
       (.I0(A1[3]),
        .I1(a11),
        .O(D[3]));
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[4]_i_1 
       (.I0(A1[4]),
        .I1(a11),
        .O(D[4]));
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[5]_i_1 
       (.I0(A1[5]),
        .I1(a11),
        .O(D[5]));
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \a1d[6]_i_1 
       (.I0(A1[6]),
        .I1(a11),
        .O(D[6]));
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a1d[7]_i_1 
       (.I0(a11),
        .I1(A1[7]),
        .O(D[7]));
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a1d[8]_i_1 
       (.I0(a11),
        .I1(A1[8]),
        .O(D[8]));
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \a1d[9]_i_1 
       (.I0(a11),
        .I1(A1[9]),
        .O(D[9]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[0] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0_n_0),
        .Q(a[0]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[10] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__9_n_0),
        .Q(a[10]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[11] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__10_n_0),
        .Q(a[11]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[1] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__0_n_0),
        .Q(a[1]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[2] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__1_n_0),
        .Q(a[2]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[3] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__2_n_0),
        .Q(a[3]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[4] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__3_n_0),
        .Q(a[4]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[5] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__4_n_0),
        .Q(a[5]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[6] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__5_n_0),
        .Q(a[6]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[7] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__6_n_0),
        .Q(a[7]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[8] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__7_n_0),
        .Q(a[8]));
  FDCE #(
    .INIT(1'b0)) 
    \a_reg[9] 
       (.C(clk_i),
        .CE(a_0),
        .CLR(rst_i),
        .D(g0_b0__8_n_0),
        .Q(a[9]));
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \b1d[0]_i_1 
       (.I0(B1[0]),
        .I1(b11),
        .O(\B1_reg[11]_0 [0]));
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \b1d[10]_i_1 
       (.I0(B1[10]),
        .I1(b11),
        .O(\B1_reg[11]_0 [10]));
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[11]_i_1 
       (.I0(b11),
        .I1(B1[11]),
        .O(\B1_reg[11]_0 [11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAABAAAA)) 
    \b1d[11]_i_2 
       (.I0(Q),
        .I1(\a0d_reg[11] [1]),
        .I2(\a0d_reg[11] [0]),
        .I3(\a0d_reg[11] [2]),
        .I4(sh[3]),
        .I5(\b1d[11]_i_3_n_0 ),
        .O(b11));
  LUT5 #(
    .INIT(32'h3E800280)) 
    \b1d[11]_i_3 
       (.I0(sh[1]),
        .I1(\a0d_reg[11] [1]),
        .I2(\a0d_reg[11] [0]),
        .I3(\a0d_reg[11] [2]),
        .I4(sh[2]),
        .O(\b1d[11]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[1]_i_1 
       (.I0(b11),
        .I1(B1[1]),
        .O(\B1_reg[11]_0 [1]));
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[2]_i_1 
       (.I0(b11),
        .I1(B1[2]),
        .O(\B1_reg[11]_0 [2]));
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[3]_i_1 
       (.I0(b11),
        .I1(B1[3]),
        .O(\B1_reg[11]_0 [3]));
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[4]_i_1 
       (.I0(b11),
        .I1(B1[4]),
        .O(\B1_reg[11]_0 [4]));
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[5]_i_1 
       (.I0(b11),
        .I1(B1[5]),
        .O(\B1_reg[11]_0 [5]));
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \b1d[6]_i_1 
       (.I0(B1[6]),
        .I1(b11),
        .O(\B1_reg[11]_0 [6]));
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[7]_i_1 
       (.I0(b11),
        .I1(B1[7]),
        .O(\B1_reg[11]_0 [7]));
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[8]_i_1 
       (.I0(b11),
        .I1(B1[8]),
        .O(\B1_reg[11]_0 [8]));
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \b1d[9]_i_1 
       (.I0(b11),
        .I1(B1[9]),
        .O(\B1_reg[11]_0 [9]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \fi[11]_i_1 
       (.I0(st_reg[3]),
        .I1(st_reg[2]),
        .I2(st_reg[1]),
        .I3(st_reg[4]),
        .I4(st_reg[0]),
        .O(esh));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[0] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[0]),
        .Q(fi[0]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[10] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[10]),
        .Q(fi[10]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[11] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[11]),
        .Q(fi[11]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[1] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[1]),
        .Q(fi[1]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[2] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[2]),
        .Q(fi[2]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[3] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[3]),
        .Q(fi[3]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[4] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[4]),
        .Q(fi[4]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[5] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[5]),
        .Q(fi[5]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[6] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[6]),
        .Q(fi[6]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[7] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[7]),
        .Q(fi[7]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[8] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[8]),
        .Q(fi[8]));
  FDCE #(
    .INIT(1'b0)) 
    \fi_reg[9] 
       (.C(clk_i),
        .CE(esh),
        .CLR(rst_i),
        .D(FREQ[9]),
        .Q(fi[9]));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[0]),
        .O(g0_b0_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__0
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[1]),
        .O(g0_b0__0_n_0));
  LUT5 #(
    .INIT(32'h0000FDE0)) 
    g0_b0__0__0
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .O(g0_b0__0__0_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__1
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[2]),
        .O(g0_b0__1_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__10
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[11]),
        .O(g0_b0__10_n_0));
  LUT5 #(
    .INIT(32'h00037298)) 
    g0_b0__11
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .O(a_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__2
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[3]),
        .O(g0_b0__2_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__3
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[4]),
        .O(g0_b0__3_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__4
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[5]),
        .O(g0_b0__4_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__5
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[6]),
        .O(g0_b0__5_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__6
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[7]),
        .O(g0_b0__6_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__7
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[8]),
        .O(g0_b0__7_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__8
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[9]),
        .O(g0_b0__8_n_0));
  LUT6 #(
    .INIT(64'h0003629800000000)) 
    g0_b0__9
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(q[10]),
        .O(g0_b0__9_n_0));
  LUT4 #(
    .INIT(16'h0EEE)) 
    i__carry__0_i_1__2
       (.I0(p_2_in),
        .I1(sr[10]),
        .I2(i__carry_i_18_n_0),
        .I3(a[10]),
        .O(p_1_in__1[10]));
  LUT4 #(
    .INIT(16'h0EEE)) 
    i__carry__0_i_2
       (.I0(p_2_in),
        .I1(sr[9]),
        .I2(i__carry_i_18_n_0),
        .I3(a[9]),
        .O(p_1_in__1[9]));
  LUT5 #(
    .INIT(32'h5555F033)) 
    i__carry__0_i_3
       (.I0(a[8]),
        .I1(fi[11]),
        .I2(sr[8]),
        .I3(i__carry_i_21_n_0),
        .I4(i__carry_i_18_n_0),
        .O(p_1_in__1[8]));
  LUT4 #(
    .INIT(16'h0DEE)) 
    i__carry__0_i_4
       (.I0(sr[11]),
        .I1(p_2_in),
        .I2(i__carry_i_18_n_0),
        .I3(a[11]),
        .O(i__carry__0_i_4_n_0));
  LUT5 #(
    .INIT(32'hA0B35FBC)) 
    i__carry__0_i_5
       (.I0(i__carry_i_18_n_0),
        .I1(sr[10]),
        .I2(a[10]),
        .I3(p_2_in),
        .I4(eb1),
        .O(i__carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h5BFC)) 
    i__carry__0_i_6
       (.I0(i__carry_i_18_n_0),
        .I1(sr[9]),
        .I2(p_2_in),
        .I3(a[9]),
        .O(i__carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h4051BFAEEAFBEAFB)) 
    i__carry__0_i_7
       (.I0(i__carry_i_18_n_0),
        .I1(i__carry_i_21_n_0),
        .I2(sr[8]),
        .I3(fi[11]),
        .I4(p_2_in),
        .I5(a[8]),
        .O(i__carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hA655A6AA)) 
    i__carry_i_10__2
       (.I0(p_1_in__1[7]),
        .I1(a[7]),
        .I2(i__carry_i_18_n_0),
        .I3(i__carry_i_21_n_0),
        .I4(st_reg[0]),
        .O(i__carry_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h51510051AE51FFAE)) 
    i__carry_i_11__4
       (.I0(i__carry_i_22_n_0),
        .I1(sr[6]),
        .I2(p_2_in),
        .I3(i__carry_i_18_n_0),
        .I4(a[6]),
        .I5(i__carry_i_33_n_0),
        .O(i__carry_i_11__4_n_0));
  LUT6 #(
    .INIT(64'h55A655A6555555A6)) 
    i__carry_i_12__0
       (.I0(p_1_in__1[5]),
        .I1(a[5]),
        .I2(p_2_in),
        .I3(ea0),
        .I4(st_reg[0]),
        .I5(i__carry_i_21_n_0),
        .O(i__carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'hAA9AAA9A5555AA9A)) 
    i__carry_i_13
       (.I0(p_1_in__1[4]),
        .I1(\shii[0]_i_1_n_0 ),
        .I2(st_reg[0]),
        .I3(i__carry_i_21_n_0),
        .I4(a[4]),
        .I5(p_2_in),
        .O(i__carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h55A6)) 
    i__carry_i_14
       (.I0(p_1_in__1[3]),
        .I1(a[3]),
        .I2(p_2_in),
        .I3(ea0),
        .O(i__carry_i_14_n_0));
  LUT3 #(
    .INIT(8'h9A)) 
    i__carry_i_15
       (.I0(p_1_in__1[2]),
        .I1(p_2_in),
        .I2(a[2]),
        .O(i__carry_i_15_n_0));
  LUT6 #(
    .INIT(64'hAA6AAA6A5555AA6A)) 
    i__carry_i_16
       (.I0(p_1_in__1[1]),
        .I1(\shii[0]_i_1_n_0 ),
        .I2(st_reg[0]),
        .I3(i__carry_i_21_n_0),
        .I4(a[1]),
        .I5(p_2_in),
        .O(i__carry_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFF1F1000001F10)) 
    i__carry_i_17
       (.I0(i__carry_i_34_n_0),
        .I1(i__carry_i_35_n_0),
        .I2(i__carry_i_33_n_0),
        .I3(sr[0]),
        .I4(i__carry_i_18_n_0),
        .I5(a[0]),
        .O(i__carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT5 #(
    .INIT(32'h01100010)) 
    i__carry_i_18
       (.I0(st_reg[1]),
        .I1(st_reg[3]),
        .I2(st_reg[2]),
        .I3(st_reg[4]),
        .I4(st_reg[0]),
        .O(i__carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT5 #(
    .INIT(32'hFFFF44F0)) 
    i__carry_i_19
       (.I0(fi[10]),
        .I1(fi[11]),
        .I2(sr[7]),
        .I3(i__carry_i_33_n_0),
        .I4(i__carry_i_18_n_0),
        .O(i__carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hAAA8A88AAAAAA88A)) 
    i__carry_i_1__2
       (.I0(a[0]),
        .I1(st_reg[3]),
        .I2(st_reg[2]),
        .I3(st_reg[1]),
        .I4(st_reg[4]),
        .I5(st_reg[0]),
        .O(i__carry_i_1__2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    i__carry_i_20
       (.I0(fi[9]),
        .I1(fi[10]),
        .I2(fi[11]),
        .I3(fi[8]),
        .O(i__carry_i_20_n_0));
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    i__carry_i_21
       (.I0(st_reg[4]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .O(i__carry_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000000FFF53)) 
    i__carry_i_22
       (.I0(fi[7]),
        .I1(fi[6]),
        .I2(fi[8]),
        .I3(\shii[0]_i_1_n_0 ),
        .I4(fi[9]),
        .I5(i__carry_i_21_n_0),
        .O(i__carry_i_22_n_0));
  LUT6 #(
    .INIT(64'h55555502555555F2)) 
    i__carry_i_23
       (.I0(fi[8]),
        .I1(fi[6]),
        .I2(fi[9]),
        .I3(fi[10]),
        .I4(fi[11]),
        .I5(fi[7]),
        .O(i__carry_i_23_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    i__carry_i_24
       (.I0(fi[5]),
        .I1(fi[8]),
        .I2(fi[11]),
        .I3(fi[10]),
        .I4(fi[9]),
        .O(i__carry_i_24_n_0));
  LUT6 #(
    .INIT(64'h555503005555F3F0)) 
    i__carry_i_25
       (.I0(fi[7]),
        .I1(fi[5]),
        .I2(fi[9]),
        .I3(fi[8]),
        .I4(\shii[0]_i_1_n_0 ),
        .I5(fi[6]),
        .O(i__carry_i_25_n_0));
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    i__carry_i_26
       (.I0(fi[4]),
        .I1(fi[8]),
        .I2(fi[11]),
        .I3(fi[10]),
        .I4(fi[9]),
        .O(i__carry_i_26_n_0));
  LUT6 #(
    .INIT(64'h555503005555F3F0)) 
    i__carry_i_27
       (.I0(fi[6]),
        .I1(fi[4]),
        .I2(fi[9]),
        .I3(fi[8]),
        .I4(\shii[0]_i_1_n_0 ),
        .I5(fi[5]),
        .O(i__carry_i_27_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    i__carry_i_28
       (.I0(fi[3]),
        .I1(fi[8]),
        .I2(fi[11]),
        .I3(fi[10]),
        .I4(fi[9]),
        .O(i__carry_i_28_n_0));
  LUT6 #(
    .INIT(64'h555503005555F3F0)) 
    i__carry_i_29
       (.I0(fi[5]),
        .I1(fi[3]),
        .I2(fi[9]),
        .I3(fi[8]),
        .I4(\shii[0]_i_1_n_0 ),
        .I5(fi[4]),
        .O(i__carry_i_29_n_0));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    i__carry_i_2__2
       (.I0(i__carry_i_18_n_0),
        .I1(a[7]),
        .I2(i__carry_i_19_n_0),
        .I3(i__carry_i_20_n_0),
        .I4(i__carry_i_21_n_0),
        .I5(fi[7]),
        .O(p_1_in__1[7]));
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    i__carry_i_30
       (.I0(fi[2]),
        .I1(fi[8]),
        .I2(fi[11]),
        .I3(fi[10]),
        .I4(fi[9]),
        .O(i__carry_i_30_n_0));
  LUT6 #(
    .INIT(64'h555503005555F3F0)) 
    i__carry_i_31
       (.I0(fi[4]),
        .I1(fi[2]),
        .I2(fi[9]),
        .I3(fi[8]),
        .I4(\shii[0]_i_1_n_0 ),
        .I5(fi[3]),
        .O(i__carry_i_31_n_0));
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    i__carry_i_32
       (.I0(fi[1]),
        .I1(fi[8]),
        .I2(fi[11]),
        .I3(fi[10]),
        .I4(fi[9]),
        .O(i__carry_i_32_n_0));
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    i__carry_i_33
       (.I0(st_reg[3]),
        .I1(st_reg[2]),
        .I2(st_reg[1]),
        .I3(st_reg[4]),
        .O(i__carry_i_33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    i__carry_i_34
       (.I0(fi[0]),
        .I1(fi[8]),
        .I2(fi[11]),
        .I3(fi[10]),
        .I4(fi[9]),
        .O(i__carry_i_34_n_0));
  LUT6 #(
    .INIT(64'h555503005555F3F0)) 
    i__carry_i_35
       (.I0(fi[3]),
        .I1(fi[1]),
        .I2(fi[9]),
        .I3(fi[8]),
        .I4(\shii[0]_i_1_n_0 ),
        .I5(fi[2]),
        .O(i__carry_i_35_n_0));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    i__carry_i_3__2
       (.I0(i__carry_i_22_n_0),
        .I1(sr[6]),
        .I2(p_2_in),
        .I3(i__carry_i_18_n_0),
        .I4(a[6]),
        .O(p_1_in__1[6]));
  LUT6 #(
    .INIT(64'h7477747774777444)) 
    i__carry_i_4__2
       (.I0(a[5]),
        .I1(i__carry_i_18_n_0),
        .I2(sr[5]),
        .I3(i__carry_i_21_n_0),
        .I4(i__carry_i_23_n_0),
        .I5(i__carry_i_24_n_0),
        .O(p_1_in__1[5]));
  LUT6 #(
    .INIT(64'h7477747774777444)) 
    i__carry_i_5__2
       (.I0(a[4]),
        .I1(i__carry_i_18_n_0),
        .I2(sr[4]),
        .I3(i__carry_i_21_n_0),
        .I4(i__carry_i_25_n_0),
        .I5(i__carry_i_26_n_0),
        .O(p_1_in__1[4]));
  LUT6 #(
    .INIT(64'h7477747774777444)) 
    i__carry_i_6__1
       (.I0(a[3]),
        .I1(i__carry_i_18_n_0),
        .I2(sr[3]),
        .I3(i__carry_i_21_n_0),
        .I4(i__carry_i_27_n_0),
        .I5(i__carry_i_28_n_0),
        .O(p_1_in__1[3]));
  LUT6 #(
    .INIT(64'h7477747774777444)) 
    i__carry_i_7__1
       (.I0(a[2]),
        .I1(i__carry_i_18_n_0),
        .I2(sr[2]),
        .I3(i__carry_i_21_n_0),
        .I4(i__carry_i_29_n_0),
        .I5(i__carry_i_30_n_0),
        .O(p_1_in__1[2]));
  LUT6 #(
    .INIT(64'h7477747774777444)) 
    i__carry_i_8__0
       (.I0(a[1]),
        .I1(i__carry_i_18_n_0),
        .I2(sr[1]),
        .I3(i__carry_i_21_n_0),
        .I4(i__carry_i_31_n_0),
        .I5(i__carry_i_32_n_0),
        .O(p_1_in__1[1]));
  LUT5 #(
    .INIT(32'h00000338)) 
    i__carry_i_9__1
       (.I0(st_reg[0]),
        .I1(st_reg[4]),
        .I2(st_reg[1]),
        .I3(st_reg[2]),
        .I4(st_reg[3]),
        .O(p_2_in));
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \shii[0]_i_1 
       (.I0(fi[10]),
        .I1(fi[11]),
        .O(\shii[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \shii[1]_i_1 
       (.I0(fi[9]),
        .I1(fi[10]),
        .I2(fi[11]),
        .O(shi[1]));
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \shii[2]_i_1 
       (.I0(fi[9]),
        .I1(fi[8]),
        .I2(fi[10]),
        .I3(fi[11]),
        .O(shi[2]));
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \shii[3]_i_1 
       (.I0(fi[8]),
        .I1(fi[11]),
        .I2(fi[10]),
        .I3(fi[9]),
        .O(shi[3]));
  FDPE #(
    .INIT(1'b1)) 
    \shii_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\shii[0]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(Q));
  FDCE #(
    .INIT(1'b0)) 
    \shii_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(shi[1]),
        .Q(sh[1]));
  FDCE #(
    .INIT(1'b0)) 
    \shii_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(shi[2]),
        .Q(sh[2]));
  FDCE #(
    .INIT(1'b0)) 
    \shii_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(shi[3]),
        .Q(sh[3]));
  LUT4 #(
    .INIT(16'h88B8)) 
    \sr[0]_i_1 
       (.I0(a[0]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[1]),
        .I3(\sr[10]_i_3_n_0 ),
        .O(\sr[0]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[10]_i_1 
       (.I0(a[10]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[9]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[11]),
        .O(\sr[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT5 #(
    .INIT(32'h00021000)) 
    \sr[10]_i_2 
       (.I0(st_reg[3]),
        .I1(st_reg[4]),
        .I2(st_reg[2]),
        .I3(st_reg[0]),
        .I4(st_reg[1]),
        .O(\sr[10]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT5 #(
    .INIT(32'h000001A0)) 
    \sr[10]_i_3 
       (.I0(st_reg[1]),
        .I1(st_reg[0]),
        .I2(st_reg[2]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .O(\sr[10]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAACFAAC0)) 
    \sr[11]_i_1 
       (.I0(a[11]),
        .I1(sr[10]),
        .I2(\sr[10]_i_3_n_0 ),
        .I3(\sr[10]_i_2_n_0 ),
        .I4(sr[11]),
        .O(\sr[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[1]_i_1 
       (.I0(a[1]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[0]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[2]),
        .O(\sr[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[2]_i_1 
       (.I0(a[2]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[1]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[3]),
        .O(\sr[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[3]_i_1 
       (.I0(a[3]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[2]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[4]),
        .O(\sr[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_1 
       (.I0(a[4]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[3]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[5]),
        .O(\sr[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[5]_i_1 
       (.I0(a[5]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[4]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[6]),
        .O(\sr[5]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[6]_i_1 
       (.I0(a[6]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[5]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[7]),
        .O(\sr[6]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[7]_i_1 
       (.I0(a[7]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[6]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[8]),
        .O(\sr[7]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[8]_i_1 
       (.I0(a[8]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[7]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[9]),
        .O(\sr[8]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[9]_i_1 
       (.I0(a[9]),
        .I1(\sr[10]_i_2_n_0 ),
        .I2(sr[8]),
        .I3(\sr[10]_i_3_n_0 ),
        .I4(sr[10]),
        .O(\sr[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[0] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[0]_i_1_n_0 ),
        .Q(sr[0]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[10] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[10]_i_1_n_0 ),
        .Q(sr[10]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\sr[11]_i_1_n_0 ),
        .Q(sr[11]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[1] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[1]_i_1_n_0 ),
        .Q(sr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[2] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[2]_i_1_n_0 ),
        .Q(sr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[3] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[3]_i_1_n_0 ),
        .Q(sr[3]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[4] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[4]_i_1_n_0 ),
        .Q(sr[4]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[5] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[5]_i_1_n_0 ),
        .Q(sr[5]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[6] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[6]_i_1_n_0 ),
        .Q(sr[6]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[7] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[7]_i_1_n_0 ),
        .Q(sr[7]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[8] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[8]_i_1_n_0 ),
        .Q(sr[8]));
  FDCE #(
    .INIT(1'b0)) 
    \sr_reg[9] 
       (.C(clk_i),
        .CE(g0_b0__0__0_n_0),
        .CLR(rst_i),
        .D(\sr[9]_i_1_n_0 ),
        .Q(sr[9]));
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \st[0]_i_1 
       (.I0(st_reg[0]),
        .O(plusOp__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \st[1]_i_1 
       (.I0(st_reg[0]),
        .I1(st_reg[1]),
        .O(plusOp__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \st[2]_i_1 
       (.I0(st_reg[1]),
        .I1(st_reg[2]),
        .I2(st_reg[0]),
        .O(plusOp__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \st[3]_i_1 
       (.I0(st_reg[3]),
        .I1(st_reg[1]),
        .I2(st_reg[2]),
        .I3(st_reg[0]),
        .O(\st[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \st[4]_i_1 
       (.I0(st_reg[0]),
        .I1(st_reg[2]),
        .I2(st_reg[1]),
        .I3(st_reg[3]),
        .I4(st_reg[4]),
        .I5(out),
        .O(\st[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \st[4]_i_2 
       (.I0(st_reg[4]),
        .I1(st_reg[0]),
        .I2(st_reg[2]),
        .I3(st_reg[1]),
        .I4(st_reg[3]),
        .O(plusOp__0[4]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[0] 
       (.C(clk_i),
        .CE(\st[4]_i_1_n_0 ),
        .CLR(rst_i),
        .D(plusOp__0[0]),
        .Q(st_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[1] 
       (.C(clk_i),
        .CE(\st[4]_i_1_n_0 ),
        .CLR(rst_i),
        .D(plusOp__0[1]),
        .Q(st_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[2] 
       (.C(clk_i),
        .CE(\st[4]_i_1_n_0 ),
        .CLR(rst_i),
        .D(plusOp__0[2]),
        .Q(st_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[3] 
       (.C(clk_i),
        .CE(\st[4]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\st[3]_i_1_n_0 ),
        .Q(st_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[4] 
       (.C(clk_i),
        .CE(\st[4]_i_1_n_0 ),
        .CLR(rst_i),
        .D(plusOp__0[4]),
        .Q(st_reg[4]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY
   (clk_i_0,
    D,
    Q,
    S,
    \z1d1_reg[15] ,
    clk_i);
  output [15:0]clk_i_0;
  output [17:0]D;
  input [19:0]Q;
  input [4:0]S;
  input [15:0]\z1d1_reg[15] ;
  input clk_i;

  wire [17:0]D;
  wire [19:0]Q;
  wire [4:0]S;
  wire clk_i;
  wire [15:0]clk_i_0;
  wire \tt2_z1[15]_i_2_n_0 ;
  wire \tt2_z1[15]_i_3_n_0 ;
  wire \tt2_z1[15]_i_4_n_0 ;
  wire \tt2_z1[15]_i_5_n_0 ;
  wire \tt2_z1[15]_i_6_n_0 ;
  wire \tt2_z1[15]_i_7_n_0 ;
  wire \tt2_z1[15]_i_8_n_0 ;
  wire \tt2_z1[15]_i_9_n_0 ;
  wire \tt2_z1[7]_i_2_n_0 ;
  wire \tt2_z1[7]_i_3_n_0 ;
  wire \tt2_z1[7]_i_4_n_0 ;
  wire \tt2_z1[7]_i_5_n_0 ;
  wire \tt2_z1[7]_i_6_n_0 ;
  wire \tt2_z1[7]_i_7_n_0 ;
  wire \tt2_z1[7]_i_8_n_0 ;
  wire \tt2_z1[7]_i_9_n_0 ;
  wire \tt2_z1_reg[15]_i_1_n_0 ;
  wire \tt2_z1_reg[15]_i_1_n_1 ;
  wire \tt2_z1_reg[15]_i_1_n_2 ;
  wire \tt2_z1_reg[15]_i_1_n_3 ;
  wire \tt2_z1_reg[15]_i_1_n_4 ;
  wire \tt2_z1_reg[15]_i_1_n_5 ;
  wire \tt2_z1_reg[15]_i_1_n_6 ;
  wire \tt2_z1_reg[15]_i_1_n_7 ;
  wire \tt2_z1_reg[21]_i_1_n_3 ;
  wire \tt2_z1_reg[21]_i_1_n_4 ;
  wire \tt2_z1_reg[21]_i_1_n_5 ;
  wire \tt2_z1_reg[21]_i_1_n_6 ;
  wire \tt2_z1_reg[21]_i_1_n_7 ;
  wire \tt2_z1_reg[7]_i_1_n_0 ;
  wire \tt2_z1_reg[7]_i_1_n_1 ;
  wire \tt2_z1_reg[7]_i_1_n_2 ;
  wire \tt2_z1_reg[7]_i_1_n_3 ;
  wire \tt2_z1_reg[7]_i_1_n_4 ;
  wire \tt2_z1_reg[7]_i_1_n_5 ;
  wire \tt2_z1_reg[7]_i_1_n_6 ;
  wire \tt2_z1_reg[7]_i_1_n_7 ;
  wire [15:0]\z1d1_reg[15] ;
  wire [7:5]\NLW_tt2_z1_reg[21]_i_1_CO_UNCONNECTED ;
  wire [7:6]\NLW_tt2_z1_reg[21]_i_1_O_UNCONNECTED ;
  wire [3:0]\NLW_tt2_z1_reg[7]_i_1_O_UNCONNECTED ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [0]),
        .Q(clk_i_0[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [10]),
        .Q(clk_i_0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [11]),
        .Q(clk_i_0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [12]),
        .Q(clk_i_0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [13]),
        .Q(clk_i_0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [14]),
        .Q(clk_i_0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [15]),
        .Q(clk_i_0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [1]),
        .Q(clk_i_0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [2]),
        .Q(clk_i_0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [3]),
        .Q(clk_i_0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [4]),
        .Q(clk_i_0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [5]),
        .Q(clk_i_0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [6]),
        .Q(clk_i_0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [7]),
        .Q(clk_i_0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [8]),
        .Q(clk_i_0[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z1d1_reg[15] [9]),
        .Q(clk_i_0[9]));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_2 
       (.I0(Q[15]),
        .I1(clk_i_0[15]),
        .O(\tt2_z1[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_3 
       (.I0(Q[14]),
        .I1(clk_i_0[14]),
        .O(\tt2_z1[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_4 
       (.I0(Q[13]),
        .I1(clk_i_0[13]),
        .O(\tt2_z1[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_5 
       (.I0(Q[12]),
        .I1(clk_i_0[12]),
        .O(\tt2_z1[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_6 
       (.I0(Q[11]),
        .I1(clk_i_0[11]),
        .O(\tt2_z1[15]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_7 
       (.I0(Q[10]),
        .I1(clk_i_0[10]),
        .O(\tt2_z1[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_8 
       (.I0(Q[9]),
        .I1(clk_i_0[9]),
        .O(\tt2_z1[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[15]_i_9 
       (.I0(Q[8]),
        .I1(clk_i_0[8]),
        .O(\tt2_z1[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_2 
       (.I0(Q[7]),
        .I1(clk_i_0[7]),
        .O(\tt2_z1[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_3 
       (.I0(Q[6]),
        .I1(clk_i_0[6]),
        .O(\tt2_z1[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_4 
       (.I0(Q[5]),
        .I1(clk_i_0[5]),
        .O(\tt2_z1[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_5 
       (.I0(Q[4]),
        .I1(clk_i_0[4]),
        .O(\tt2_z1[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_6 
       (.I0(Q[3]),
        .I1(clk_i_0[3]),
        .O(\tt2_z1[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_7 
       (.I0(Q[2]),
        .I1(clk_i_0[2]),
        .O(\tt2_z1[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_8 
       (.I0(Q[1]),
        .I1(clk_i_0[1]),
        .O(\tt2_z1[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2_z1[7]_i_9 
       (.I0(Q[0]),
        .I1(clk_i_0[0]),
        .O(\tt2_z1[7]_i_9_n_0 ));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tt2_z1_reg[15]_i_1 
       (.CI(\tt2_z1_reg[7]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tt2_z1_reg[15]_i_1_n_0 ,\tt2_z1_reg[15]_i_1_n_1 ,\tt2_z1_reg[15]_i_1_n_2 ,\tt2_z1_reg[15]_i_1_n_3 ,\tt2_z1_reg[15]_i_1_n_4 ,\tt2_z1_reg[15]_i_1_n_5 ,\tt2_z1_reg[15]_i_1_n_6 ,\tt2_z1_reg[15]_i_1_n_7 }),
        .DI(Q[15:8]),
        .O(D[11:4]),
        .S({\tt2_z1[15]_i_2_n_0 ,\tt2_z1[15]_i_3_n_0 ,\tt2_z1[15]_i_4_n_0 ,\tt2_z1[15]_i_5_n_0 ,\tt2_z1[15]_i_6_n_0 ,\tt2_z1[15]_i_7_n_0 ,\tt2_z1[15]_i_8_n_0 ,\tt2_z1[15]_i_9_n_0 }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tt2_z1_reg[21]_i_1 
       (.CI(\tt2_z1_reg[15]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_tt2_z1_reg[21]_i_1_CO_UNCONNECTED [7:5],\tt2_z1_reg[21]_i_1_n_3 ,\tt2_z1_reg[21]_i_1_n_4 ,\tt2_z1_reg[21]_i_1_n_5 ,\tt2_z1_reg[21]_i_1_n_6 ,\tt2_z1_reg[21]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,Q[19:16]}),
        .O({\NLW_tt2_z1_reg[21]_i_1_O_UNCONNECTED [7:6],D[17:12]}),
        .S({1'b0,1'b0,1'b1,S}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tt2_z1_reg[7]_i_1 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\tt2_z1_reg[7]_i_1_n_0 ,\tt2_z1_reg[7]_i_1_n_1 ,\tt2_z1_reg[7]_i_1_n_2 ,\tt2_z1_reg[7]_i_1_n_3 ,\tt2_z1_reg[7]_i_1_n_4 ,\tt2_z1_reg[7]_i_1_n_5 ,\tt2_z1_reg[7]_i_1_n_6 ,\tt2_z1_reg[7]_i_1_n_7 }),
        .DI(Q[7:0]),
        .O({D[3:0],\NLW_tt2_z1_reg[7]_i_1_O_UNCONNECTED [3:0]}),
        .S({\tt2_z1[7]_i_2_n_0 ,\tt2_z1[7]_i_3_n_0 ,\tt2_z1[7]_i_4_n_0 ,\tt2_z1[7]_i_5_n_0 ,\tt2_z1[7]_i_6_n_0 ,\tt2_z1[7]_i_7_n_0 ,\tt2_z1[7]_i_8_n_0 ,\tt2_z1[7]_i_9_n_0 }));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY_0
   (Q,
    SE11_out,
    D,
    clk_i);
  output [15:0]Q;
  input SE11_out;
  input [15:0]D;
  input clk_i;

  wire [15:0]D;
  wire [15:0]Q;
  wire SE11_out;
  wire clk_i;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[0]),
        .Q(Q[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[10]),
        .Q(Q[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[11]),
        .Q(Q[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[12]),
        .Q(Q[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[13]),
        .Q(Q[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[14]),
        .Q(Q[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[15]),
        .Q(Q[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[1]),
        .Q(Q[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[2]),
        .Q(Q[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[3]),
        .Q(Q[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[4]),
        .Q(Q[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[5]),
        .Q(Q[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[6]),
        .Q(Q[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[7]),
        .Q(Q[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[8]),
        .Q(Q[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_56/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[9]),
        .Q(Q[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized1
   (Q,
    SE11_out,
    D,
    clk_i);
  output [15:0]Q;
  input SE11_out;
  input [15:0]D;
  input clk_i;

  wire [15:0]D;
  wire [15:0]Q;
  wire SE11_out;
  wire clk_i;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[0]),
        .Q(Q[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[10]),
        .Q(Q[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[11]),
        .Q(Q[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[12]),
        .Q(Q[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[13]),
        .Q(Q[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[14]),
        .Q(Q[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[15]),
        .Q(Q[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[1]),
        .Q(Q[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[2]),
        .Q(Q[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[3]),
        .Q(Q[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[4]),
        .Q(Q[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[5]),
        .Q(Q[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[6]),
        .Q(Q[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[7]),
        .Q(Q[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[8]),
        .Q(Q[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_56/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[9]),
        .Q(Q[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized11
   (SE,
    D,
    clk_i_0,
    Q,
    P,
    \d3_3_reg[15] ,
    clk_i);
  output SE;
  output [15:0]D;
  output [15:0]clk_i_0;
  input [1:0]Q;
  input [15:0]P;
  input [15:0]\d3_3_reg[15] ;
  input clk_i;

  wire [15:0]D;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_1 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_2 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_3 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_4 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_5 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_6 ;
  wire \D16.DEL0[0].U_SRL_i_1__5_n_7 ;
  wire \D16.DEL0[0].U_SRL_i_2__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_3__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_4__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_5__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_6__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_7__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_8__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_9__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_1 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_2 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_3 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_4 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_5 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_6 ;
  wire \D16.DEL0[8].U_SRL_i_1__3_n_7 ;
  wire \D16.DEL0[8].U_SRL_i_2_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_3_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_4_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_5_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_6_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_7_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_8_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_9_n_0 ;
  wire [15:0]P;
  wire [1:0]Q;
  wire SE;
  wire clk_i;
  wire [15:0]clk_i_0;
  wire [15:0]\d3_3_reg[15] ;
  wire [7:7]\NLW_D16.DEL0[8].U_SRL_i_1__3_CO_UNCONNECTED ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[0]),
        .Q(clk_i_0[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \D16.DEL0[0].U_SRL_i_1__1 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(SE));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[0].U_SRL_i_1__5 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\D16.DEL0[0].U_SRL_i_1__5_n_0 ,\D16.DEL0[0].U_SRL_i_1__5_n_1 ,\D16.DEL0[0].U_SRL_i_1__5_n_2 ,\D16.DEL0[0].U_SRL_i_1__5_n_3 ,\D16.DEL0[0].U_SRL_i_1__5_n_4 ,\D16.DEL0[0].U_SRL_i_1__5_n_5 ,\D16.DEL0[0].U_SRL_i_1__5_n_6 ,\D16.DEL0[0].U_SRL_i_1__5_n_7 }),
        .DI(P[7:0]),
        .O(D[7:0]),
        .S({\D16.DEL0[0].U_SRL_i_2__2_n_0 ,\D16.DEL0[0].U_SRL_i_3__1_n_0 ,\D16.DEL0[0].U_SRL_i_4__0_n_0 ,\D16.DEL0[0].U_SRL_i_5__0_n_0 ,\D16.DEL0[0].U_SRL_i_6__0_n_0 ,\D16.DEL0[0].U_SRL_i_7__0_n_0 ,\D16.DEL0[0].U_SRL_i_8__0_n_0 ,\D16.DEL0[0].U_SRL_i_9__0_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_2__2 
       (.I0(P[7]),
        .I1(\d3_3_reg[15] [7]),
        .O(\D16.DEL0[0].U_SRL_i_2__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_3__1 
       (.I0(P[6]),
        .I1(\d3_3_reg[15] [6]),
        .O(\D16.DEL0[0].U_SRL_i_3__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_4__0 
       (.I0(P[5]),
        .I1(\d3_3_reg[15] [5]),
        .O(\D16.DEL0[0].U_SRL_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_5__0 
       (.I0(P[4]),
        .I1(\d3_3_reg[15] [4]),
        .O(\D16.DEL0[0].U_SRL_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_6__0 
       (.I0(P[3]),
        .I1(\d3_3_reg[15] [3]),
        .O(\D16.DEL0[0].U_SRL_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_7__0 
       (.I0(P[2]),
        .I1(\d3_3_reg[15] [2]),
        .O(\D16.DEL0[0].U_SRL_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_8__0 
       (.I0(P[1]),
        .I1(\d3_3_reg[15] [1]),
        .O(\D16.DEL0[0].U_SRL_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_9__0 
       (.I0(P[0]),
        .I1(\d3_3_reg[15] [0]),
        .O(\D16.DEL0[0].U_SRL_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[10]),
        .Q(clk_i_0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[11]),
        .Q(clk_i_0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[12]),
        .Q(clk_i_0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[13]),
        .Q(clk_i_0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[14]),
        .Q(clk_i_0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[15]),
        .Q(clk_i_0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[1]),
        .Q(clk_i_0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[2]),
        .Q(clk_i_0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[3]),
        .Q(clk_i_0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[4]),
        .Q(clk_i_0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[5]),
        .Q(clk_i_0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[6]),
        .Q(clk_i_0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[7]),
        .Q(clk_i_0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[8]),
        .Q(clk_i_0[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[8].U_SRL_i_1__3 
       (.CI(\D16.DEL0[0].U_SRL_i_1__5_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_D16.DEL0[8].U_SRL_i_1__3_CO_UNCONNECTED [7],\D16.DEL0[8].U_SRL_i_1__3_n_1 ,\D16.DEL0[8].U_SRL_i_1__3_n_2 ,\D16.DEL0[8].U_SRL_i_1__3_n_3 ,\D16.DEL0[8].U_SRL_i_1__3_n_4 ,\D16.DEL0[8].U_SRL_i_1__3_n_5 ,\D16.DEL0[8].U_SRL_i_1__3_n_6 ,\D16.DEL0[8].U_SRL_i_1__3_n_7 }),
        .DI({1'b0,P[14:8]}),
        .O(D[15:8]),
        .S({\D16.DEL0[8].U_SRL_i_2_n_0 ,\D16.DEL0[8].U_SRL_i_3_n_0 ,\D16.DEL0[8].U_SRL_i_4_n_0 ,\D16.DEL0[8].U_SRL_i_5_n_0 ,\D16.DEL0[8].U_SRL_i_6_n_0 ,\D16.DEL0[8].U_SRL_i_7_n_0 ,\D16.DEL0[8].U_SRL_i_8_n_0 ,\D16.DEL0[8].U_SRL_i_9_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_2 
       (.I0(P[15]),
        .I1(\d3_3_reg[15] [15]),
        .O(\D16.DEL0[8].U_SRL_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_3 
       (.I0(P[14]),
        .I1(\d3_3_reg[15] [14]),
        .O(\D16.DEL0[8].U_SRL_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_4 
       (.I0(P[13]),
        .I1(\d3_3_reg[15] [13]),
        .O(\D16.DEL0[8].U_SRL_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_5 
       (.I0(P[12]),
        .I1(\d3_3_reg[15] [12]),
        .O(\D16.DEL0[8].U_SRL_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_6 
       (.I0(P[11]),
        .I1(\d3_3_reg[15] [11]),
        .O(\D16.DEL0[8].U_SRL_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_7 
       (.I0(P[10]),
        .I1(\d3_3_reg[15] [10]),
        .O(\D16.DEL0[8].U_SRL_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_8 
       (.I0(P[9]),
        .I1(\d3_3_reg[15] [9]),
        .O(\D16.DEL0[8].U_SRL_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_9 
       (.I0(P[8]),
        .I1(\d3_3_reg[15] [8]),
        .O(\D16.DEL0[8].U_SRL_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_78/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[9]),
        .Q(clk_i_0[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized13
   (D,
    Q,
    \D32.DEL1[15].U_SRL0_0 ,
    \D32.DEL1[15].U_SRL0_1 ,
    d4_4,
    \D32.DEL1[0].U_SRL0_0 ,
    \D32.DEL1[1].U_SRL0_0 ,
    \D32.DEL1[2].U_SRL0_0 ,
    \D32.DEL1[3].U_SRL0_0 ,
    \D32.DEL1[4].U_SRL0_0 ,
    \D32.DEL1[5].U_SRL0_0 ,
    \D32.DEL1[6].U_SRL0_0 ,
    \D32.DEL1[7].U_SRL0_0 ,
    \D32.DEL1[8].U_SRL0_0 ,
    \D32.DEL1[9].U_SRL0_0 ,
    \D32.DEL1[10].U_SRL0_0 ,
    \D32.DEL1[11].U_SRL0_0 ,
    \D32.DEL1[12].U_SRL0_0 ,
    \D32.DEL1[13].U_SRL0_0 ,
    \D32.DEL1[14].U_SRL0_0 ,
    \D32.DEL1[15].U_SRL0_2 ,
    \D32.DEL1[15].U_SRL1_0 ,
    clk_i);
  output [15:0]D;
  input [2:0]Q;
  input \D32.DEL1[15].U_SRL0_0 ;
  input \D32.DEL1[15].U_SRL0_1 ;
  input [15:0]d4_4;
  input \D32.DEL1[0].U_SRL0_0 ;
  input \D32.DEL1[1].U_SRL0_0 ;
  input \D32.DEL1[2].U_SRL0_0 ;
  input \D32.DEL1[3].U_SRL0_0 ;
  input \D32.DEL1[4].U_SRL0_0 ;
  input \D32.DEL1[5].U_SRL0_0 ;
  input \D32.DEL1[6].U_SRL0_0 ;
  input \D32.DEL1[7].U_SRL0_0 ;
  input \D32.DEL1[8].U_SRL0_0 ;
  input \D32.DEL1[9].U_SRL0_0 ;
  input \D32.DEL1[10].U_SRL0_0 ;
  input \D32.DEL1[11].U_SRL0_0 ;
  input \D32.DEL1[12].U_SRL0_0 ;
  input \D32.DEL1[13].U_SRL0_0 ;
  input \D32.DEL1[14].U_SRL0_0 ;
  input \D32.DEL1[15].U_SRL0_2 ;
  input [15:0]\D32.DEL1[15].U_SRL1_0 ;
  input clk_i;

  wire [15:0]D;
  wire \D32.DEL1[0].U_SRL0_0 ;
  wire \D32.DEL1[10].U_SRL0_0 ;
  wire \D32.DEL1[11].U_SRL0_0 ;
  wire \D32.DEL1[12].U_SRL0_0 ;
  wire \D32.DEL1[13].U_SRL0_0 ;
  wire \D32.DEL1[14].U_SRL0_0 ;
  wire \D32.DEL1[15].U_SRL0_0 ;
  wire \D32.DEL1[15].U_SRL0_1 ;
  wire \D32.DEL1[15].U_SRL0_2 ;
  wire [15:0]\D32.DEL1[15].U_SRL1_0 ;
  wire \D32.DEL1[1].U_SRL0_0 ;
  wire \D32.DEL1[2].U_SRL0_0 ;
  wire \D32.DEL1[3].U_SRL0_0 ;
  wire \D32.DEL1[4].U_SRL0_0 ;
  wire \D32.DEL1[5].U_SRL0_0 ;
  wire \D32.DEL1[6].U_SRL0_0 ;
  wire \D32.DEL1[7].U_SRL0_0 ;
  wire \D32.DEL1[8].U_SRL0_0 ;
  wire \D32.DEL1[9].U_SRL0_0 ;
  wire [2:0]Q;
  wire SE2_out;
  wire clk_i;
  wire [15:0]d4_4;
  wire [15:0]d78_4;
  wire di1_0;
  wire di1_1;
  wire di1_10;
  wire di1_11;
  wire di1_12;
  wire di1_13;
  wire di1_14;
  wire di1_15;
  wire di1_2;
  wire di1_3;
  wire di1_4;
  wire di1_5;
  wire di1_6;
  wire di1_7;
  wire di1_8;
  wire di1_9;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[0].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[0].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [0]),
        .Q(di1_0));
  LUT3 #(
    .INIT(8'h06)) 
    \D32.DEL1[0].U_SRL0_i_1 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .O(SE2_out));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[0].U_SRL0_i_1__0 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[0]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[0]),
        .I4(\D32.DEL1[0].U_SRL0_0 ),
        .O(D[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[0].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[0].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_0),
        .Q(d78_4[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[10].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[10].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [10]),
        .Q(di1_10));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[10].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[10]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[10]),
        .I4(\D32.DEL1[10].U_SRL0_0 ),
        .O(D[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[10].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[10].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_10),
        .Q(d78_4[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[11].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[11].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [11]),
        .Q(di1_11));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[11].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[11]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[11]),
        .I4(\D32.DEL1[11].U_SRL0_0 ),
        .O(D[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[11].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[11].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_11),
        .Q(d78_4[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[12].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[12].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [12]),
        .Q(di1_12));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[12].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[12]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[12]),
        .I4(\D32.DEL1[12].U_SRL0_0 ),
        .O(D[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[12].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[12].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_12),
        .Q(d78_4[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[13].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[13].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [13]),
        .Q(di1_13));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[13].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[13]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[13]),
        .I4(\D32.DEL1[13].U_SRL0_0 ),
        .O(D[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[13].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[13].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_13),
        .Q(d78_4[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[14].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[14].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [14]),
        .Q(di1_14));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[14].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[14]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[14]),
        .I4(\D32.DEL1[14].U_SRL0_0 ),
        .O(D[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[14].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[14].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_14),
        .Q(d78_4[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[15].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[15].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [15]),
        .Q(di1_15));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[15].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[15]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[15]),
        .I4(\D32.DEL1[15].U_SRL0_2 ),
        .O(D[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[15].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[15].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_15),
        .Q(d78_4[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[1].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[1].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [1]),
        .Q(di1_1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[1].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[1]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[1]),
        .I4(\D32.DEL1[1].U_SRL0_0 ),
        .O(D[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[1].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[1].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_1),
        .Q(d78_4[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[2].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[2].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [2]),
        .Q(di1_2));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[2].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[2]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[2]),
        .I4(\D32.DEL1[2].U_SRL0_0 ),
        .O(D[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[2].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[2].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_2),
        .Q(d78_4[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[3].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[3].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [3]),
        .Q(di1_3));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[3].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[3]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[3]),
        .I4(\D32.DEL1[3].U_SRL0_0 ),
        .O(D[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[3].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[3].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_3),
        .Q(d78_4[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[4].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[4].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [4]),
        .Q(di1_4));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[4].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[4]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[4]),
        .I4(\D32.DEL1[4].U_SRL0_0 ),
        .O(D[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[4].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[4].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_4),
        .Q(d78_4[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[5].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[5].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [5]),
        .Q(di1_5));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[5].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[5]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[5]),
        .I4(\D32.DEL1[5].U_SRL0_0 ),
        .O(D[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[5].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[5].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_5),
        .Q(d78_4[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[6].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[6].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [6]),
        .Q(di1_6));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[6].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[6]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[6]),
        .I4(\D32.DEL1[6].U_SRL0_0 ),
        .O(D[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[6].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[6].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_6),
        .Q(d78_4[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[7].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[7].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [7]),
        .Q(di1_7));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[7].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[7]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[7]),
        .I4(\D32.DEL1[7].U_SRL0_0 ),
        .O(D[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[7].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[7].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_7),
        .Q(d78_4[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[8].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[8].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [8]),
        .Q(di1_8));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[8].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[8]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[8]),
        .I4(\D32.DEL1[8].U_SRL0_0 ),
        .O(D[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[8].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[8].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_8),
        .Q(d78_4[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[9].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[9].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL1_0 [9]),
        .Q(di1_9));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \D32.DEL1[9].U_SRL0_i_1 
       (.I0(\D32.DEL1[15].U_SRL0_0 ),
        .I1(d78_4[9]),
        .I2(\D32.DEL1[15].U_SRL0_1 ),
        .I3(d4_4[9]),
        .I4(\D32.DEL1[9].U_SRL0_0 ),
        .O(D[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_78/D32.DEL1[9].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[9].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(SE2_out),
        .CLK(clk_i),
        .D(di1_9),
        .Q(d78_4[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized16
   (Q,
    D,
    clk_i);
  output [15:0]Q;
  input [15:0]D;
  input clk_i;

  wire [15:0]D;
  wire [15:0]Q;
  wire clk_i;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[0]),
        .Q(Q[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[10]),
        .Q(Q[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[11]),
        .Q(Q[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[12]),
        .Q(Q[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[13]),
        .Q(Q[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[14]),
        .Q(Q[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[15]),
        .Q(Q[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[1]),
        .Q(Q[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[2]),
        .Q(Q[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[3]),
        .Q(Q[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[4]),
        .Q(Q[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[5]),
        .Q(Q[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[6]),
        .Q(Q[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[7]),
        .Q(Q[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[8]),
        .Q(Q[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[9]),
        .Q(Q[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized18
   (clk_i_0,
    O,
    \st_reg[2] ,
    doii1,
    Q,
    \DO_reg[15] ,
    D,
    clk_i);
  output [15:0]clk_i_0;
  output [1:0]O;
  output \st_reg[2] ;
  input doii1;
  input [2:0]Q;
  input [18:0]\DO_reg[15] ;
  input [15:0]D;
  input clk_i;

  wire [15:0]D;
  wire \D16.DEL0[0].U_SRL_i_10_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_11_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_1 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_2 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_3 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_4 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_5 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_6 ;
  wire \D16.DEL0[0].U_SRL_i_3__0_n_7 ;
  wire \D16.DEL0[0].U_SRL_i_4_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_5_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_6_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_7_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_8_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_9_n_0 ;
  wire \D16.DEL0[15].U_SRL_i_2_n_6 ;
  wire \D16.DEL0[15].U_SRL_i_2_n_7 ;
  wire \D16.DEL0[7].U_SRL_i_10_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_1 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_2 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_3 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_4 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_5 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_6 ;
  wire \D16.DEL0[7].U_SRL_i_2_n_7 ;
  wire \D16.DEL0[7].U_SRL_i_3_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_4_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_5_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_6_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_7_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_8_n_0 ;
  wire \D16.DEL0[7].U_SRL_i_9_n_0 ;
  wire [18:0]\DO_reg[15] ;
  wire [1:0]O;
  wire [2:0]Q;
  wire clk_i;
  wire [15:0]clk_i_0;
  wire di1_0;
  wire di1_1;
  wire di1_10;
  wire di1_11;
  wire di1_12;
  wire di1_13;
  wire di1_14;
  wire di1_15;
  wire di1_2;
  wire di1_3;
  wire di1_4;
  wire di1_5;
  wire di1_6;
  wire di1_7;
  wire di1_8;
  wire di1_9;
  wire doii1;
  wire [16:1]plusOp18;
  wire \st_reg[2] ;
  wire [15:0]z4;
  wire [0:0]\NLW_D16.DEL0[0].U_SRL_i_3__0_O_UNCONNECTED ;
  wire [7:2]\NLW_D16.DEL0[15].U_SRL_i_2_CO_UNCONNECTED ;
  wire [7:3]\NLW_D16.DEL0[15].U_SRL_i_2_O_UNCONNECTED ;

  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_10 
       (.I0(z4[1]),
        .I1(\DO_reg[15] [1]),
        .O(\D16.DEL0[0].U_SRL_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_11 
       (.I0(z4[0]),
        .I1(\DO_reg[15] [0]),
        .O(\D16.DEL0[0].U_SRL_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[0].U_SRL_i_1__0 
       (.I0(z4[0]),
        .I1(doii1),
        .I2(plusOp18[1]),
        .O(clk_i_0[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[0].U_SRL_i_3__0 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\D16.DEL0[0].U_SRL_i_3__0_n_0 ,\D16.DEL0[0].U_SRL_i_3__0_n_1 ,\D16.DEL0[0].U_SRL_i_3__0_n_2 ,\D16.DEL0[0].U_SRL_i_3__0_n_3 ,\D16.DEL0[0].U_SRL_i_3__0_n_4 ,\D16.DEL0[0].U_SRL_i_3__0_n_5 ,\D16.DEL0[0].U_SRL_i_3__0_n_6 ,\D16.DEL0[0].U_SRL_i_3__0_n_7 }),
        .DI(z4[7:0]),
        .O({plusOp18[7:1],\NLW_D16.DEL0[0].U_SRL_i_3__0_O_UNCONNECTED [0]}),
        .S({\D16.DEL0[0].U_SRL_i_4_n_0 ,\D16.DEL0[0].U_SRL_i_5_n_0 ,\D16.DEL0[0].U_SRL_i_6_n_0 ,\D16.DEL0[0].U_SRL_i_7_n_0 ,\D16.DEL0[0].U_SRL_i_8_n_0 ,\D16.DEL0[0].U_SRL_i_9_n_0 ,\D16.DEL0[0].U_SRL_i_10_n_0 ,\D16.DEL0[0].U_SRL_i_11_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_4 
       (.I0(z4[7]),
        .I1(\DO_reg[15] [7]),
        .O(\D16.DEL0[0].U_SRL_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_5 
       (.I0(z4[6]),
        .I1(\DO_reg[15] [6]),
        .O(\D16.DEL0[0].U_SRL_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_6 
       (.I0(z4[5]),
        .I1(\DO_reg[15] [5]),
        .O(\D16.DEL0[0].U_SRL_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_7 
       (.I0(z4[4]),
        .I1(\DO_reg[15] [4]),
        .O(\D16.DEL0[0].U_SRL_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_8 
       (.I0(z4[3]),
        .I1(\DO_reg[15] [3]),
        .O(\D16.DEL0[0].U_SRL_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_9 
       (.I0(z4[2]),
        .I1(\DO_reg[15] [2]),
        .O(\D16.DEL0[0].U_SRL_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[10].U_SRL_i_1 
       (.I0(z4[10]),
        .I1(doii1),
        .I2(plusOp18[11]),
        .O(clk_i_0[10]));
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[11].U_SRL_i_1 
       (.I0(z4[11]),
        .I1(doii1),
        .I2(plusOp18[12]),
        .O(clk_i_0[11]));
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[12].U_SRL_i_1 
       (.I0(z4[12]),
        .I1(doii1),
        .I2(plusOp18[13]),
        .O(clk_i_0[12]));
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[13].U_SRL_i_1 
       (.I0(z4[13]),
        .I1(doii1),
        .I2(plusOp18[14]),
        .O(clk_i_0[13]));
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[14].U_SRL_i_1 
       (.I0(z4[14]),
        .I1(doii1),
        .I2(plusOp18[15]),
        .O(clk_i_0[14]));
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[15].U_SRL_i_1 
       (.I0(z4[15]),
        .I1(doii1),
        .I2(plusOp18[16]),
        .O(clk_i_0[15]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[15].U_SRL_i_2 
       (.CI(\D16.DEL0[7].U_SRL_i_2_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_D16.DEL0[15].U_SRL_i_2_CO_UNCONNECTED [7:2],\D16.DEL0[15].U_SRL_i_2_n_6 ,\D16.DEL0[15].U_SRL_i_2_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_D16.DEL0[15].U_SRL_i_2_O_UNCONNECTED [7:3],O,plusOp18[16]}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,\DO_reg[15] [18:16]}));
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[1].U_SRL_i_1 
       (.I0(z4[1]),
        .I1(doii1),
        .I2(plusOp18[2]),
        .O(clk_i_0[1]));
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[2].U_SRL_i_1 
       (.I0(z4[2]),
        .I1(doii1),
        .I2(plusOp18[3]),
        .O(clk_i_0[2]));
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[3].U_SRL_i_1 
       (.I0(z4[3]),
        .I1(doii1),
        .I2(plusOp18[4]),
        .O(clk_i_0[3]));
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[4].U_SRL_i_1 
       (.I0(z4[4]),
        .I1(doii1),
        .I2(plusOp18[5]),
        .O(clk_i_0[4]));
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[5].U_SRL_i_1 
       (.I0(z4[5]),
        .I1(doii1),
        .I2(plusOp18[6]),
        .O(clk_i_0[5]));
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[6].U_SRL_i_1 
       (.I0(z4[6]),
        .I1(doii1),
        .I2(plusOp18[7]),
        .O(clk_i_0[6]));
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[7].U_SRL_i_1 
       (.I0(z4[7]),
        .I1(doii1),
        .I2(plusOp18[8]),
        .O(clk_i_0[7]));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_10 
       (.I0(z4[8]),
        .I1(\DO_reg[15] [8]),
        .O(\D16.DEL0[7].U_SRL_i_10_n_0 ));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[7].U_SRL_i_2 
       (.CI(\D16.DEL0[0].U_SRL_i_3__0_n_0 ),
        .CI_TOP(1'b0),
        .CO({\D16.DEL0[7].U_SRL_i_2_n_0 ,\D16.DEL0[7].U_SRL_i_2_n_1 ,\D16.DEL0[7].U_SRL_i_2_n_2 ,\D16.DEL0[7].U_SRL_i_2_n_3 ,\D16.DEL0[7].U_SRL_i_2_n_4 ,\D16.DEL0[7].U_SRL_i_2_n_5 ,\D16.DEL0[7].U_SRL_i_2_n_6 ,\D16.DEL0[7].U_SRL_i_2_n_7 }),
        .DI(z4[15:8]),
        .O(plusOp18[15:8]),
        .S({\D16.DEL0[7].U_SRL_i_3_n_0 ,\D16.DEL0[7].U_SRL_i_4_n_0 ,\D16.DEL0[7].U_SRL_i_5_n_0 ,\D16.DEL0[7].U_SRL_i_6_n_0 ,\D16.DEL0[7].U_SRL_i_7_n_0 ,\D16.DEL0[7].U_SRL_i_8_n_0 ,\D16.DEL0[7].U_SRL_i_9_n_0 ,\D16.DEL0[7].U_SRL_i_10_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_3 
       (.I0(z4[15]),
        .I1(\DO_reg[15] [15]),
        .O(\D16.DEL0[7].U_SRL_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_4 
       (.I0(z4[14]),
        .I1(\DO_reg[15] [14]),
        .O(\D16.DEL0[7].U_SRL_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_5 
       (.I0(z4[13]),
        .I1(\DO_reg[15] [13]),
        .O(\D16.DEL0[7].U_SRL_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_6 
       (.I0(z4[12]),
        .I1(\DO_reg[15] [12]),
        .O(\D16.DEL0[7].U_SRL_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_7 
       (.I0(z4[11]),
        .I1(\DO_reg[15] [11]),
        .O(\D16.DEL0[7].U_SRL_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_8 
       (.I0(z4[10]),
        .I1(\DO_reg[15] [10]),
        .O(\D16.DEL0[7].U_SRL_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[7].U_SRL_i_9 
       (.I0(z4[9]),
        .I1(\DO_reg[15] [9]),
        .O(\D16.DEL0[7].U_SRL_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[8].U_SRL_i_1 
       (.I0(z4[8]),
        .I1(doii1),
        .I2(plusOp18[9]),
        .O(clk_i_0[8]));
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D16.DEL0[9].U_SRL_i_1 
       (.I0(z4[9]),
        .I1(doii1),
        .I2(plusOp18[10]),
        .O(clk_i_0[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[0].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[0].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[0]),
        .Q(di1_0));
  LUT3 #(
    .INIT(8'h14)) 
    \D32.DEL1[0].U_SRL0_i_2 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\st_reg[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[0].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[0].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_0),
        .Q(z4[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[10].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[10].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[10]),
        .Q(di1_10));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[10].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[10].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_10),
        .Q(z4[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[11].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[11].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[11]),
        .Q(di1_11));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[11].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[11].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_11),
        .Q(z4[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[12].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[12].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[12]),
        .Q(di1_12));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[12].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[12].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_12),
        .Q(z4[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[13].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[13].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[13]),
        .Q(di1_13));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[13].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[13].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_13),
        .Q(z4[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[14].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[14].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[14]),
        .Q(di1_14));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[14].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[14].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_14),
        .Q(z4[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[15].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[15].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[15]),
        .Q(di1_15));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[15].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[15].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_15),
        .Q(z4[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[1].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[1].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[1]),
        .Q(di1_1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[1].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[1].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_1),
        .Q(z4[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[2].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[2].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[2]),
        .Q(di1_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[2].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[2].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_2),
        .Q(z4[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[3].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[3].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[3]),
        .Q(di1_3));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[3].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[3].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_3),
        .Q(z4[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[4].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[4].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[4]),
        .Q(di1_4));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[4].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[4].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_4),
        .Q(z4[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[5].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[5].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[5]),
        .Q(di1_5));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[5].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[5].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_5),
        .Q(z4[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[6].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[6].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[6]),
        .Q(di1_6));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[6].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[6].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_6),
        .Q(z4[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[7].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[7].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[7]),
        .Q(di1_7));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[7].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[7].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_7),
        .Q(z4[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[8].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[8].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[8]),
        .Q(di1_8));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[8].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[8].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_8),
        .Q(z4[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[9].U_SRL0 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[9].U_SRL0 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b1),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(D[9]),
        .Q(di1_9));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4/D32.DEL1[9].U_SRL1 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D32.DEL1[9].U_SRL1 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(di1_9),
        .Q(z4[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized20
   (D,
    \did_reg[15] ,
    Q,
    \d_z2_reg[15] ,
    \dd1_reg[15] ,
    DI,
    S,
    \dd1_reg[15]_0 ,
    clk_i);
  output [15:0]D;
  output [16:0]\did_reg[15] ;
  input [2:0]Q;
  input [15:0]\d_z2_reg[15] ;
  input [13:0]\dd1_reg[15] ;
  input [1:0]DI;
  input [2:0]S;
  input [15:0]\dd1_reg[15]_0 ;
  input clk_i;

  wire [15:0]D;
  wire \D16.DEL0[0].U_SRL_n_0 ;
  wire \D16.DEL0[10].U_SRL_n_0 ;
  wire \D16.DEL0[11].U_SRL_n_0 ;
  wire \D16.DEL0[12].U_SRL_n_0 ;
  wire \D16.DEL0[13].U_SRL_n_0 ;
  wire \D16.DEL0[14].U_SRL_n_0 ;
  wire \D16.DEL0[15].U_SRL_n_0 ;
  wire \D16.DEL0[1].U_SRL_n_0 ;
  wire \D16.DEL0[2].U_SRL_n_0 ;
  wire \D16.DEL0[3].U_SRL_n_0 ;
  wire \D16.DEL0[4].U_SRL_n_0 ;
  wire \D16.DEL0[5].U_SRL_n_0 ;
  wire \D16.DEL0[6].U_SRL_n_0 ;
  wire \D16.DEL0[7].U_SRL_n_0 ;
  wire \D16.DEL0[8].U_SRL_n_0 ;
  wire \D16.DEL0[9].U_SRL_n_0 ;
  wire [1:0]DI;
  wire [2:0]Q;
  wire [2:0]S;
  wire clk_i;
  wire \d_z2[15]_i_2_n_0 ;
  wire \d_z2[15]_i_3_n_0 ;
  wire \d_z2[15]_i_4_n_0 ;
  wire \d_z2[15]_i_5_n_0 ;
  wire \d_z2[15]_i_6_n_0 ;
  wire \d_z2[15]_i_7_n_0 ;
  wire \d_z2[15]_i_8_n_0 ;
  wire \d_z2[15]_i_9_n_0 ;
  wire \d_z2[7]_i_10_n_0 ;
  wire \d_z2[7]_i_11_n_0 ;
  wire \d_z2[7]_i_2_n_0 ;
  wire \d_z2[7]_i_3_n_0 ;
  wire \d_z2[7]_i_4_n_0 ;
  wire \d_z2[7]_i_5_n_0 ;
  wire \d_z2[7]_i_6_n_0 ;
  wire \d_z2[7]_i_7_n_0 ;
  wire \d_z2[7]_i_8_n_0 ;
  wire \d_z2[7]_i_9_n_0 ;
  wire [15:0]\d_z2_reg[15] ;
  wire \d_z2_reg[15]_i_1_n_0 ;
  wire \d_z2_reg[15]_i_1_n_1 ;
  wire \d_z2_reg[15]_i_1_n_2 ;
  wire \d_z2_reg[15]_i_1_n_3 ;
  wire \d_z2_reg[15]_i_1_n_4 ;
  wire \d_z2_reg[15]_i_1_n_5 ;
  wire \d_z2_reg[15]_i_1_n_6 ;
  wire \d_z2_reg[15]_i_1_n_7 ;
  wire \d_z2_reg[20]_i_1_n_5 ;
  wire \d_z2_reg[20]_i_1_n_6 ;
  wire \d_z2_reg[20]_i_1_n_7 ;
  wire \d_z2_reg[7]_i_1_n_0 ;
  wire \d_z2_reg[7]_i_1_n_1 ;
  wire \d_z2_reg[7]_i_1_n_2 ;
  wire \d_z2_reg[7]_i_1_n_3 ;
  wire \d_z2_reg[7]_i_1_n_4 ;
  wire \d_z2_reg[7]_i_1_n_5 ;
  wire \d_z2_reg[7]_i_1_n_6 ;
  wire \d_z2_reg[7]_i_1_n_7 ;
  wire [13:0]\dd1_reg[15] ;
  wire [15:0]\dd1_reg[15]_0 ;
  wire [16:0]\did_reg[15] ;
  wire [7:3]\NLW_d_z2_reg[20]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_d_z2_reg[20]_i_1_O_UNCONNECTED ;
  wire [2:0]\NLW_d_z2_reg[7]_i_1_O_UNCONNECTED ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [0]),
        .Q(\D16.DEL0[0].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [10]),
        .Q(\D16.DEL0[10].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [11]),
        .Q(\D16.DEL0[11].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [12]),
        .Q(\D16.DEL0[12].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [13]),
        .Q(\D16.DEL0[13].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [14]),
        .Q(\D16.DEL0[14].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [15]),
        .Q(\D16.DEL0[15].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [1]),
        .Q(\D16.DEL0[1].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [2]),
        .Q(\D16.DEL0[2].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [3]),
        .Q(\D16.DEL0[3].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [4]),
        .Q(\D16.DEL0[4].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [5]),
        .Q(\D16.DEL0[5].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [6]),
        .Q(\D16.DEL0[6].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [7]),
        .Q(\D16.DEL0[7].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [8]),
        .Q(\D16.DEL0[8].U_SRL_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DD/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DD/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b0),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\dd1_reg[15]_0 [9]),
        .Q(\D16.DEL0[9].U_SRL_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_2 
       (.I0(\D16.DEL0[15].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [13]),
        .I5(\d_z2_reg[15] [15]),
        .O(\d_z2[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_3 
       (.I0(\D16.DEL0[14].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [12]),
        .I5(\d_z2_reg[15] [14]),
        .O(\d_z2[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_4 
       (.I0(\D16.DEL0[13].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [11]),
        .I5(\d_z2_reg[15] [13]),
        .O(\d_z2[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_5 
       (.I0(\D16.DEL0[12].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [10]),
        .I5(\d_z2_reg[15] [12]),
        .O(\d_z2[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_6 
       (.I0(\D16.DEL0[11].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [9]),
        .I5(\d_z2_reg[15] [11]),
        .O(\d_z2[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_7 
       (.I0(\D16.DEL0[10].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [8]),
        .I5(\d_z2_reg[15] [10]),
        .O(\d_z2[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_8 
       (.I0(\D16.DEL0[9].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [7]),
        .I5(\d_z2_reg[15] [9]),
        .O(\d_z2[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[15]_i_9 
       (.I0(\D16.DEL0[8].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [6]),
        .I5(\d_z2_reg[15] [8]),
        .O(\d_z2[15]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFD0002FF)) 
    \d_z2[7]_i_10 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(\D16.DEL0[1].U_SRL_n_0 ),
        .I4(\d_z2_reg[15] [1]),
        .O(\d_z2[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFD0002FF)) 
    \d_z2[7]_i_11 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(\D16.DEL0[0].U_SRL_n_0 ),
        .I4(\d_z2_reg[15] [0]),
        .O(\d_z2[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \d_z2[7]_i_2 
       (.I0(\D16.DEL0[1].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\d_z2[7]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \d_z2[7]_i_3 
       (.I0(\D16.DEL0[0].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\d_z2[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[7]_i_4 
       (.I0(\D16.DEL0[7].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [5]),
        .I5(\d_z2_reg[15] [7]),
        .O(\d_z2[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[7]_i_5 
       (.I0(\D16.DEL0[6].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [4]),
        .I5(\d_z2_reg[15] [6]),
        .O(\d_z2[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[7]_i_6 
       (.I0(\D16.DEL0[5].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [3]),
        .I5(\d_z2_reg[15] [5]),
        .O(\d_z2[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[7]_i_7 
       (.I0(\D16.DEL0[4].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [2]),
        .I5(\d_z2_reg[15] [4]),
        .O(\d_z2[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[7]_i_8 
       (.I0(\D16.DEL0[3].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [1]),
        .I5(\d_z2_reg[15] [3]),
        .O(\d_z2[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hABAAA8AA54555755)) 
    \d_z2[7]_i_9 
       (.I0(\D16.DEL0[2].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\dd1_reg[15] [0]),
        .I5(\d_z2_reg[15] [2]),
        .O(\d_z2[7]_i_9_n_0 ));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \d_z2_reg[15]_i_1 
       (.CI(\d_z2_reg[7]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\d_z2_reg[15]_i_1_n_0 ,\d_z2_reg[15]_i_1_n_1 ,\d_z2_reg[15]_i_1_n_2 ,\d_z2_reg[15]_i_1_n_3 ,\d_z2_reg[15]_i_1_n_4 ,\d_z2_reg[15]_i_1_n_5 ,\d_z2_reg[15]_i_1_n_6 ,\d_z2_reg[15]_i_1_n_7 }),
        .DI(D[15:8]),
        .O(\did_reg[15] [12:5]),
        .S({\d_z2[15]_i_2_n_0 ,\d_z2[15]_i_3_n_0 ,\d_z2[15]_i_4_n_0 ,\d_z2[15]_i_5_n_0 ,\d_z2[15]_i_6_n_0 ,\d_z2[15]_i_7_n_0 ,\d_z2[15]_i_8_n_0 ,\d_z2[15]_i_9_n_0 }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \d_z2_reg[20]_i_1 
       (.CI(\d_z2_reg[15]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_d_z2_reg[20]_i_1_CO_UNCONNECTED [7:3],\d_z2_reg[20]_i_1_n_5 ,\d_z2_reg[20]_i_1_n_6 ,\d_z2_reg[20]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,DI}),
        .O({\NLW_d_z2_reg[20]_i_1_O_UNCONNECTED [7:4],\did_reg[15] [16:13]}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b1,S}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \d_z2_reg[7]_i_1 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\d_z2_reg[7]_i_1_n_0 ,\d_z2_reg[7]_i_1_n_1 ,\d_z2_reg[7]_i_1_n_2 ,\d_z2_reg[7]_i_1_n_3 ,\d_z2_reg[7]_i_1_n_4 ,\d_z2_reg[7]_i_1_n_5 ,\d_z2_reg[7]_i_1_n_6 ,\d_z2_reg[7]_i_1_n_7 }),
        .DI({D[7:2],\d_z2[7]_i_2_n_0 ,\d_z2[7]_i_3_n_0 }),
        .O({\did_reg[15] [4:0],\NLW_d_z2_reg[7]_i_1_O_UNCONNECTED [2:0]}),
        .S({\d_z2[7]_i_4_n_0 ,\d_z2[7]_i_5_n_0 ,\d_z2[7]_i_6_n_0 ,\d_z2[7]_i_7_n_0 ,\d_z2[7]_i_8_n_0 ,\d_z2[7]_i_9_n_0 ,\d_z2[7]_i_10_n_0 ,\d_z2[7]_i_11_n_0 }));
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT4 #(
    .INIT(16'hA8AA)) 
    \dd1[0]_i_1 
       (.I0(\D16.DEL0[0].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(D[0]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[10]_i_1 
       (.I0(\dd1_reg[15] [8]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[10].U_SRL_n_0 ),
        .O(D[10]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[11]_i_1 
       (.I0(\dd1_reg[15] [9]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[11].U_SRL_n_0 ),
        .O(D[11]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[12]_i_1 
       (.I0(\dd1_reg[15] [10]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[12].U_SRL_n_0 ),
        .O(D[12]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[13]_i_1 
       (.I0(\dd1_reg[15] [11]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[13].U_SRL_n_0 ),
        .O(D[13]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[14]_i_1 
       (.I0(\dd1_reg[15] [12]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[14].U_SRL_n_0 ),
        .O(D[14]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[15]_i_1 
       (.I0(\dd1_reg[15] [13]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[15].U_SRL_n_0 ),
        .O(D[15]));
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT4 #(
    .INIT(16'hA8AA)) 
    \dd1[1]_i_1 
       (.I0(\D16.DEL0[1].U_SRL_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(D[1]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[2]_i_1 
       (.I0(\dd1_reg[15] [0]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[2].U_SRL_n_0 ),
        .O(D[2]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[3]_i_1 
       (.I0(\dd1_reg[15] [1]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[3].U_SRL_n_0 ),
        .O(D[3]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[4]_i_1 
       (.I0(\dd1_reg[15] [2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[4].U_SRL_n_0 ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[5]_i_1 
       (.I0(\dd1_reg[15] [3]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[5].U_SRL_n_0 ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[6]_i_1 
       (.I0(\dd1_reg[15] [4]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[6].U_SRL_n_0 ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[7]_i_1 
       (.I0(\dd1_reg[15] [5]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[7].U_SRL_n_0 ),
        .O(D[7]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[8]_i_1 
       (.I0(\dd1_reg[15] [6]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[8].U_SRL_n_0 ),
        .O(D[8]));
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \dd1[9]_i_1 
       (.I0(\dd1_reg[15] [7]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(\D16.DEL0[9].U_SRL_n_0 ),
        .O(D[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized3
   (clk_i_0,
    D,
    Q,
    S,
    \z3d1_reg[15] ,
    clk_i);
  output [15:0]clk_i_0;
  output [17:0]D;
  input [18:0]Q;
  input [3:0]S;
  input [15:0]\z3d1_reg[15] ;
  input clk_i;

  wire [17:0]D;
  wire [18:0]Q;
  wire [3:0]S;
  wire clk_i;
  wire [15:0]clk_i_0;
  wire \t2z2_z3[15]_i_2_n_0 ;
  wire \t2z2_z3[15]_i_3_n_0 ;
  wire \t2z2_z3[15]_i_4_n_0 ;
  wire \t2z2_z3[15]_i_5_n_0 ;
  wire \t2z2_z3[15]_i_6_n_0 ;
  wire \t2z2_z3[15]_i_7_n_0 ;
  wire \t2z2_z3[15]_i_8_n_0 ;
  wire \t2z2_z3[15]_i_9_n_0 ;
  wire \t2z2_z3[7]_i_2_n_0 ;
  wire \t2z2_z3[7]_i_3_n_0 ;
  wire \t2z2_z3[7]_i_4_n_0 ;
  wire \t2z2_z3[7]_i_5_n_0 ;
  wire \t2z2_z3[7]_i_6_n_0 ;
  wire \t2z2_z3[7]_i_7_n_0 ;
  wire \t2z2_z3[7]_i_8_n_0 ;
  wire \t2z2_z3[7]_i_9_n_0 ;
  wire \t2z2_z3_reg[15]_i_1_n_0 ;
  wire \t2z2_z3_reg[15]_i_1_n_1 ;
  wire \t2z2_z3_reg[15]_i_1_n_2 ;
  wire \t2z2_z3_reg[15]_i_1_n_3 ;
  wire \t2z2_z3_reg[15]_i_1_n_4 ;
  wire \t2z2_z3_reg[15]_i_1_n_5 ;
  wire \t2z2_z3_reg[15]_i_1_n_6 ;
  wire \t2z2_z3_reg[15]_i_1_n_7 ;
  wire \t2z2_z3_reg[19]_i_1_n_5 ;
  wire \t2z2_z3_reg[19]_i_1_n_6 ;
  wire \t2z2_z3_reg[19]_i_1_n_7 ;
  wire \t2z2_z3_reg[7]_i_1_n_0 ;
  wire \t2z2_z3_reg[7]_i_1_n_1 ;
  wire \t2z2_z3_reg[7]_i_1_n_2 ;
  wire \t2z2_z3_reg[7]_i_1_n_3 ;
  wire \t2z2_z3_reg[7]_i_1_n_4 ;
  wire \t2z2_z3_reg[7]_i_1_n_5 ;
  wire \t2z2_z3_reg[7]_i_1_n_6 ;
  wire \t2z2_z3_reg[7]_i_1_n_7 ;
  wire [15:0]\z3d1_reg[15] ;
  wire [7:3]\NLW_t2z2_z3_reg[19]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_t2z2_z3_reg[19]_i_1_O_UNCONNECTED ;
  wire [1:0]\NLW_t2z2_z3_reg[7]_i_1_O_UNCONNECTED ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [0]),
        .Q(clk_i_0[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [10]),
        .Q(clk_i_0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [11]),
        .Q(clk_i_0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [12]),
        .Q(clk_i_0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [13]),
        .Q(clk_i_0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [14]),
        .Q(clk_i_0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [15]),
        .Q(clk_i_0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [1]),
        .Q(clk_i_0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [2]),
        .Q(clk_i_0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [3]),
        .Q(clk_i_0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [4]),
        .Q(clk_i_0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [5]),
        .Q(clk_i_0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [6]),
        .Q(clk_i_0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [7]),
        .Q(clk_i_0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [8]),
        .Q(clk_i_0[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(\z3d1_reg[15] [9]),
        .Q(clk_i_0[9]));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_2 
       (.I0(Q[15]),
        .I1(clk_i_0[15]),
        .O(\t2z2_z3[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_3 
       (.I0(Q[14]),
        .I1(clk_i_0[14]),
        .O(\t2z2_z3[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_4 
       (.I0(Q[13]),
        .I1(clk_i_0[13]),
        .O(\t2z2_z3[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_5 
       (.I0(Q[12]),
        .I1(clk_i_0[12]),
        .O(\t2z2_z3[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_6 
       (.I0(Q[11]),
        .I1(clk_i_0[11]),
        .O(\t2z2_z3[15]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_7 
       (.I0(Q[10]),
        .I1(clk_i_0[10]),
        .O(\t2z2_z3[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_8 
       (.I0(Q[9]),
        .I1(clk_i_0[9]),
        .O(\t2z2_z3[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[15]_i_9 
       (.I0(Q[8]),
        .I1(clk_i_0[8]),
        .O(\t2z2_z3[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_2 
       (.I0(Q[7]),
        .I1(clk_i_0[7]),
        .O(\t2z2_z3[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_3 
       (.I0(Q[6]),
        .I1(clk_i_0[6]),
        .O(\t2z2_z3[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_4 
       (.I0(Q[5]),
        .I1(clk_i_0[5]),
        .O(\t2z2_z3[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_5 
       (.I0(Q[4]),
        .I1(clk_i_0[4]),
        .O(\t2z2_z3[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_6 
       (.I0(Q[3]),
        .I1(clk_i_0[3]),
        .O(\t2z2_z3[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_7 
       (.I0(Q[2]),
        .I1(clk_i_0[2]),
        .O(\t2z2_z3[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_8 
       (.I0(Q[1]),
        .I1(clk_i_0[1]),
        .O(\t2z2_z3[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \t2z2_z3[7]_i_9 
       (.I0(Q[0]),
        .I1(clk_i_0[0]),
        .O(\t2z2_z3[7]_i_9_n_0 ));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t2z2_z3_reg[15]_i_1 
       (.CI(\t2z2_z3_reg[7]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\t2z2_z3_reg[15]_i_1_n_0 ,\t2z2_z3_reg[15]_i_1_n_1 ,\t2z2_z3_reg[15]_i_1_n_2 ,\t2z2_z3_reg[15]_i_1_n_3 ,\t2z2_z3_reg[15]_i_1_n_4 ,\t2z2_z3_reg[15]_i_1_n_5 ,\t2z2_z3_reg[15]_i_1_n_6 ,\t2z2_z3_reg[15]_i_1_n_7 }),
        .DI(Q[15:8]),
        .O(D[13:6]),
        .S({\t2z2_z3[15]_i_2_n_0 ,\t2z2_z3[15]_i_3_n_0 ,\t2z2_z3[15]_i_4_n_0 ,\t2z2_z3[15]_i_5_n_0 ,\t2z2_z3[15]_i_6_n_0 ,\t2z2_z3[15]_i_7_n_0 ,\t2z2_z3[15]_i_8_n_0 ,\t2z2_z3[15]_i_9_n_0 }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t2z2_z3_reg[19]_i_1 
       (.CI(\t2z2_z3_reg[15]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_t2z2_z3_reg[19]_i_1_CO_UNCONNECTED [7:3],\t2z2_z3_reg[19]_i_1_n_5 ,\t2z2_z3_reg[19]_i_1_n_6 ,\t2z2_z3_reg[19]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,Q[18:16]}),
        .O({\NLW_t2z2_z3_reg[19]_i_1_O_UNCONNECTED [7:4],D[17:14]}),
        .S({1'b0,1'b0,1'b0,1'b0,S}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t2z2_z3_reg[7]_i_1 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\t2z2_z3_reg[7]_i_1_n_0 ,\t2z2_z3_reg[7]_i_1_n_1 ,\t2z2_z3_reg[7]_i_1_n_2 ,\t2z2_z3_reg[7]_i_1_n_3 ,\t2z2_z3_reg[7]_i_1_n_4 ,\t2z2_z3_reg[7]_i_1_n_5 ,\t2z2_z3_reg[7]_i_1_n_6 ,\t2z2_z3_reg[7]_i_1_n_7 }),
        .DI(Q[7:0]),
        .O({D[5:0],\NLW_t2z2_z3_reg[7]_i_1_O_UNCONNECTED [1:0]}),
        .S({\t2z2_z3[7]_i_2_n_0 ,\t2z2_z3[7]_i_3_n_0 ,\t2z2_z3[7]_i_4_n_0 ,\t2z2_z3[7]_i_5_n_0 ,\t2z2_z3[7]_i_6_n_0 ,\t2z2_z3[7]_i_7_n_0 ,\t2z2_z3[7]_i_8_n_0 ,\t2z2_z3[7]_i_9_n_0 }));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized3_1
   (SE11_out,
    clk_i_0,
    Q,
    D,
    clk_i);
  output SE11_out;
  output [15:0]clk_i_0;
  input [1:0]Q;
  input [15:0]D;
  input clk_i;

  wire [15:0]D;
  wire [1:0]Q;
  wire SE11_out;
  wire clk_i;
  wire [15:0]clk_i_0;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[0]),
        .Q(clk_i_0[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \D16.DEL0[0].U_SRL_i_1 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(SE11_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[10]),
        .Q(clk_i_0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[11]),
        .Q(clk_i_0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[12]),
        .Q(clk_i_0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[13]),
        .Q(clk_i_0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[14]),
        .Q(clk_i_0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[15]),
        .Q(clk_i_0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[1]),
        .Q(clk_i_0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[2]),
        .Q(clk_i_0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[3]),
        .Q(clk_i_0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[4]),
        .Q(clk_i_0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[5]),
        .Q(clk_i_0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[6]),
        .Q(clk_i_0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[7]),
        .Q(clk_i_0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[8]),
        .Q(clk_i_0[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ3_56/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b0),
        .CE(SE11_out),
        .CLK(clk_i),
        .D(D[9]),
        .Q(clk_i_0[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized5
   (\dd2_reg[0] ,
    \dd2_reg[1] ,
    \dd2_reg[2] ,
    \dd2_reg[3] ,
    \dd2_reg[4] ,
    \dd2_reg[5] ,
    \dd2_reg[6] ,
    \dd2_reg[7] ,
    \dd2_reg[8] ,
    \dd2_reg[9] ,
    \dd2_reg[10] ,
    \dd2_reg[11] ,
    \dd2_reg[12] ,
    \dd2_reg[13] ,
    \dd2_reg[14] ,
    \dd2_reg[15] ,
    Q,
    \D32.DEL1[15].U_SRL0_i_1 ,
    \D32.DEL1[15].U_SRL0_i_1_0 ,
    clk_i);
  output \dd2_reg[0] ;
  output \dd2_reg[1] ;
  output \dd2_reg[2] ;
  output \dd2_reg[3] ;
  output \dd2_reg[4] ;
  output \dd2_reg[5] ;
  output \dd2_reg[6] ;
  output \dd2_reg[7] ;
  output \dd2_reg[8] ;
  output \dd2_reg[9] ;
  output \dd2_reg[10] ;
  output \dd2_reg[11] ;
  output \dd2_reg[12] ;
  output \dd2_reg[13] ;
  output \dd2_reg[14] ;
  output \dd2_reg[15] ;
  input [2:0]Q;
  input [15:0]\D32.DEL1[15].U_SRL0_i_1 ;
  input [0:0]\D32.DEL1[15].U_SRL0_i_1_0 ;
  input clk_i;

  wire \D16.DEL0[0].U_SRL_i_1__7_n_0 ;
  wire [15:0]\D32.DEL1[15].U_SRL0_i_1 ;
  wire [0:0]\D32.DEL1[15].U_SRL0_i_1_0 ;
  wire [2:0]Q;
  wire clk_i;
  wire [15:0]d56_4;
  wire \dd2_reg[0] ;
  wire \dd2_reg[10] ;
  wire \dd2_reg[11] ;
  wire \dd2_reg[12] ;
  wire \dd2_reg[13] ;
  wire \dd2_reg[14] ;
  wire \dd2_reg[15] ;
  wire \dd2_reg[1] ;
  wire \dd2_reg[2] ;
  wire \dd2_reg[3] ;
  wire \dd2_reg[4] ;
  wire \dd2_reg[5] ;
  wire \dd2_reg[6] ;
  wire \dd2_reg[7] ;
  wire \dd2_reg[8] ;
  wire \dd2_reg[9] ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [0]),
        .Q(d56_4[0]));
  LUT3 #(
    .INIT(8'h81)) 
    \D16.DEL0[0].U_SRL_i_1__7 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\D16.DEL0[0].U_SRL_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [10]),
        .Q(d56_4[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [11]),
        .Q(d56_4[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [12]),
        .Q(d56_4[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [13]),
        .Q(d56_4[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [14]),
        .Q(d56_4[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [15]),
        .Q(d56_4[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [1]),
        .Q(d56_4[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [2]),
        .Q(d56_4[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [3]),
        .Q(d56_4[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [4]),
        .Q(d56_4[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [5]),
        .Q(d56_4[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [6]),
        .Q(d56_4[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [7]),
        .Q(d56_4[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [8]),
        .Q(d56_4[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ4_56/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b1),
        .A2(1'b0),
        .A3(1'b1),
        .CE(\D16.DEL0[0].U_SRL_i_1__7_n_0 ),
        .CLK(clk_i),
        .D(\D32.DEL1[15].U_SRL0_i_1 [9]),
        .Q(d56_4[9]));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[0].U_SRL0_i_4 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [0]),
        .I1(d56_4[0]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[0] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[10].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [10]),
        .I1(d56_4[10]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[10] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[11].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [11]),
        .I1(d56_4[11]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[11] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[12].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [12]),
        .I1(d56_4[12]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[12] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[13].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [13]),
        .I1(d56_4[13]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[13] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[14].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [14]),
        .I1(d56_4[14]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[14] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[15].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [15]),
        .I1(d56_4[15]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[15] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[1].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [1]),
        .I1(d56_4[1]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[1] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[2].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [2]),
        .I1(d56_4[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[2] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[3].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [3]),
        .I1(d56_4[3]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[3] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[4].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [4]),
        .I1(d56_4[4]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[4] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[5].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [5]),
        .I1(d56_4[5]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[5] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[6].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [6]),
        .I1(d56_4[6]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[6] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[7].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [7]),
        .I1(d56_4[7]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[7] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[8].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [8]),
        .I1(d56_4[8]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[8] ));
  LUT6 #(
    .INIT(64'hCAAAA00CC00AA00C)) 
    \D32.DEL1[9].U_SRL0_i_2 
       (.I0(\D32.DEL1[15].U_SRL0_i_1 [9]),
        .I1(d56_4[9]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(\D32.DEL1[15].U_SRL0_i_1_0 ),
        .O(\dd2_reg[9] ));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized7
   (D,
    clk_i_0,
    Q,
    P,
    SE,
    clk_i);
  output [15:0]D;
  output [15:0]clk_i_0;
  input [15:0]Q;
  input [15:0]P;
  input SE;
  input clk_i;

  wire [15:0]D;
  wire \D16.DEL0[0].U_SRL_i_10__0_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_1 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_2 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_3 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_4 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_5 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_6 ;
  wire \D16.DEL0[0].U_SRL_i_2__1_n_7 ;
  wire \D16.DEL0[0].U_SRL_i_3__3_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_4__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_5__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_6__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_7__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_8__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_9__2_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_1 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_2 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_3 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_4 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_5 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_6 ;
  wire \D16.DEL0[8].U_SRL_i_1__5_n_7 ;
  wire \D16.DEL0[8].U_SRL_i_2__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_3__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_4__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_5__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_6__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_7__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_8__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_9__1_n_0 ;
  wire [15:0]P;
  wire [15:0]Q;
  wire SE;
  wire clk_i;
  wire [15:0]clk_i_0;
  wire [7:7]\NLW_D16.DEL0[8].U_SRL_i_1__5_CO_UNCONNECTED ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[0]),
        .Q(clk_i_0[0]));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_10__0 
       (.I0(Q[0]),
        .I1(P[0]),
        .O(\D16.DEL0[0].U_SRL_i_10__0_n_0 ));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[0].U_SRL_i_2__1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\D16.DEL0[0].U_SRL_i_2__1_n_0 ,\D16.DEL0[0].U_SRL_i_2__1_n_1 ,\D16.DEL0[0].U_SRL_i_2__1_n_2 ,\D16.DEL0[0].U_SRL_i_2__1_n_3 ,\D16.DEL0[0].U_SRL_i_2__1_n_4 ,\D16.DEL0[0].U_SRL_i_2__1_n_5 ,\D16.DEL0[0].U_SRL_i_2__1_n_6 ,\D16.DEL0[0].U_SRL_i_2__1_n_7 }),
        .DI(Q[7:0]),
        .O(D[7:0]),
        .S({\D16.DEL0[0].U_SRL_i_3__3_n_0 ,\D16.DEL0[0].U_SRL_i_4__2_n_0 ,\D16.DEL0[0].U_SRL_i_5__2_n_0 ,\D16.DEL0[0].U_SRL_i_6__2_n_0 ,\D16.DEL0[0].U_SRL_i_7__2_n_0 ,\D16.DEL0[0].U_SRL_i_8__2_n_0 ,\D16.DEL0[0].U_SRL_i_9__2_n_0 ,\D16.DEL0[0].U_SRL_i_10__0_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_3__3 
       (.I0(Q[7]),
        .I1(P[7]),
        .O(\D16.DEL0[0].U_SRL_i_3__3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_4__2 
       (.I0(Q[6]),
        .I1(P[6]),
        .O(\D16.DEL0[0].U_SRL_i_4__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_5__2 
       (.I0(Q[5]),
        .I1(P[5]),
        .O(\D16.DEL0[0].U_SRL_i_5__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_6__2 
       (.I0(Q[4]),
        .I1(P[4]),
        .O(\D16.DEL0[0].U_SRL_i_6__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_7__2 
       (.I0(Q[3]),
        .I1(P[3]),
        .O(\D16.DEL0[0].U_SRL_i_7__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_8__2 
       (.I0(Q[2]),
        .I1(P[2]),
        .O(\D16.DEL0[0].U_SRL_i_8__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_9__2 
       (.I0(Q[1]),
        .I1(P[1]),
        .O(\D16.DEL0[0].U_SRL_i_9__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[10]),
        .Q(clk_i_0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[11]),
        .Q(clk_i_0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[12]),
        .Q(clk_i_0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[13]),
        .Q(clk_i_0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[14]),
        .Q(clk_i_0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[15]),
        .Q(clk_i_0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[1]),
        .Q(clk_i_0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[2]),
        .Q(clk_i_0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[3]),
        .Q(clk_i_0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[4]),
        .Q(clk_i_0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[5]),
        .Q(clk_i_0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[6]),
        .Q(clk_i_0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[7]),
        .Q(clk_i_0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[8]),
        .Q(clk_i_0[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[8].U_SRL_i_1__5 
       (.CI(\D16.DEL0[0].U_SRL_i_2__1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_D16.DEL0[8].U_SRL_i_1__5_CO_UNCONNECTED [7],\D16.DEL0[8].U_SRL_i_1__5_n_1 ,\D16.DEL0[8].U_SRL_i_1__5_n_2 ,\D16.DEL0[8].U_SRL_i_1__5_n_3 ,\D16.DEL0[8].U_SRL_i_1__5_n_4 ,\D16.DEL0[8].U_SRL_i_1__5_n_5 ,\D16.DEL0[8].U_SRL_i_1__5_n_6 ,\D16.DEL0[8].U_SRL_i_1__5_n_7 }),
        .DI({1'b0,Q[14:8]}),
        .O(D[15:8]),
        .S({\D16.DEL0[8].U_SRL_i_2__1_n_0 ,\D16.DEL0[8].U_SRL_i_3__1_n_0 ,\D16.DEL0[8].U_SRL_i_4__1_n_0 ,\D16.DEL0[8].U_SRL_i_5__1_n_0 ,\D16.DEL0[8].U_SRL_i_6__1_n_0 ,\D16.DEL0[8].U_SRL_i_7__1_n_0 ,\D16.DEL0[8].U_SRL_i_8__1_n_0 ,\D16.DEL0[8].U_SRL_i_9__1_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_2__1 
       (.I0(Q[15]),
        .I1(P[15]),
        .O(\D16.DEL0[8].U_SRL_i_2__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_3__1 
       (.I0(Q[14]),
        .I1(P[14]),
        .O(\D16.DEL0[8].U_SRL_i_3__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_4__1 
       (.I0(Q[13]),
        .I1(P[13]),
        .O(\D16.DEL0[8].U_SRL_i_4__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_5__1 
       (.I0(Q[12]),
        .I1(P[12]),
        .O(\D16.DEL0[8].U_SRL_i_5__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_6__1 
       (.I0(Q[11]),
        .I1(P[11]),
        .O(\D16.DEL0[8].U_SRL_i_6__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_7__1 
       (.I0(Q[10]),
        .I1(P[10]),
        .O(\D16.DEL0[8].U_SRL_i_7__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_8__1 
       (.I0(Q[9]),
        .I1(P[9]),
        .O(\D16.DEL0[8].U_SRL_i_8__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_9__1 
       (.I0(Q[8]),
        .I1(P[8]),
        .O(\D16.DEL0[8].U_SRL_i_9__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ1_78/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[9]),
        .Q(clk_i_0[9]));
endmodule

(* ORIG_REF_NAME = "DELAY" *) 
module switch_elements_DELAY__parameterized9
   (D,
    clk_i_0,
    Q,
    P,
    SE,
    clk_i);
  output [15:0]D;
  output [15:0]clk_i_0;
  input [15:0]Q;
  input [15:0]P;
  input SE;
  input clk_i;

  wire [15:0]D;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_1 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_2 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_3 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_4 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_5 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_6 ;
  wire \D16.DEL0[0].U_SRL_i_1__6_n_7 ;
  wire \D16.DEL0[0].U_SRL_i_2__3_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_3__2_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_4__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_5__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_6__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_7__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_8__1_n_0 ;
  wire \D16.DEL0[0].U_SRL_i_9__1_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_1 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_2 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_3 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_4 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_5 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_6 ;
  wire \D16.DEL0[8].U_SRL_i_1__4_n_7 ;
  wire \D16.DEL0[8].U_SRL_i_2__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_3__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_4__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_5__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_6__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_7__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_8__0_n_0 ;
  wire \D16.DEL0[8].U_SRL_i_9__0_n_0 ;
  wire [15:0]P;
  wire [15:0]Q;
  wire SE;
  wire clk_i;
  wire [15:0]clk_i_0;
  wire [7:7]\NLW_D16.DEL0[8].U_SRL_i_1__4_CO_UNCONNECTED ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[0].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[0].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[0]),
        .Q(clk_i_0[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[0].U_SRL_i_1__6 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\D16.DEL0[0].U_SRL_i_1__6_n_0 ,\D16.DEL0[0].U_SRL_i_1__6_n_1 ,\D16.DEL0[0].U_SRL_i_1__6_n_2 ,\D16.DEL0[0].U_SRL_i_1__6_n_3 ,\D16.DEL0[0].U_SRL_i_1__6_n_4 ,\D16.DEL0[0].U_SRL_i_1__6_n_5 ,\D16.DEL0[0].U_SRL_i_1__6_n_6 ,\D16.DEL0[0].U_SRL_i_1__6_n_7 }),
        .DI(Q[7:0]),
        .O(D[7:0]),
        .S({\D16.DEL0[0].U_SRL_i_2__3_n_0 ,\D16.DEL0[0].U_SRL_i_3__2_n_0 ,\D16.DEL0[0].U_SRL_i_4__1_n_0 ,\D16.DEL0[0].U_SRL_i_5__1_n_0 ,\D16.DEL0[0].U_SRL_i_6__1_n_0 ,\D16.DEL0[0].U_SRL_i_7__1_n_0 ,\D16.DEL0[0].U_SRL_i_8__1_n_0 ,\D16.DEL0[0].U_SRL_i_9__1_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_2__3 
       (.I0(Q[7]),
        .I1(P[7]),
        .O(\D16.DEL0[0].U_SRL_i_2__3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_3__2 
       (.I0(Q[6]),
        .I1(P[6]),
        .O(\D16.DEL0[0].U_SRL_i_3__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_4__1 
       (.I0(Q[5]),
        .I1(P[5]),
        .O(\D16.DEL0[0].U_SRL_i_4__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_5__1 
       (.I0(Q[4]),
        .I1(P[4]),
        .O(\D16.DEL0[0].U_SRL_i_5__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_6__1 
       (.I0(Q[3]),
        .I1(P[3]),
        .O(\D16.DEL0[0].U_SRL_i_6__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_7__1 
       (.I0(Q[2]),
        .I1(P[2]),
        .O(\D16.DEL0[0].U_SRL_i_7__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_8__1 
       (.I0(Q[1]),
        .I1(P[1]),
        .O(\D16.DEL0[0].U_SRL_i_8__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[0].U_SRL_i_9__1 
       (.I0(Q[0]),
        .I1(P[0]),
        .O(\D16.DEL0[0].U_SRL_i_9__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[10].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[10].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[10]),
        .Q(clk_i_0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[11].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[11].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[11]),
        .Q(clk_i_0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[12].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[12].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[12]),
        .Q(clk_i_0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[13].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[13].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[13]),
        .Q(clk_i_0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[14].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[14].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[14]),
        .Q(clk_i_0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[15].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[15].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[15]),
        .Q(clk_i_0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[1].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[1].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[1]),
        .Q(clk_i_0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[2].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[2].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[2]),
        .Q(clk_i_0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[3].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[3].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[3]),
        .Q(clk_i_0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[4].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[4].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[4]),
        .Q(clk_i_0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[5].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[5].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[5]),
        .Q(clk_i_0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[6].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[6].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[6]),
        .Q(clk_i_0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[7].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[7].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[7]),
        .Q(clk_i_0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[8].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[8].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[8]),
        .Q(clk_i_0[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \D16.DEL0[8].U_SRL_i_1__4 
       (.CI(\D16.DEL0[0].U_SRL_i_1__6_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_D16.DEL0[8].U_SRL_i_1__4_CO_UNCONNECTED [7],\D16.DEL0[8].U_SRL_i_1__4_n_1 ,\D16.DEL0[8].U_SRL_i_1__4_n_2 ,\D16.DEL0[8].U_SRL_i_1__4_n_3 ,\D16.DEL0[8].U_SRL_i_1__4_n_4 ,\D16.DEL0[8].U_SRL_i_1__4_n_5 ,\D16.DEL0[8].U_SRL_i_1__4_n_6 ,\D16.DEL0[8].U_SRL_i_1__4_n_7 }),
        .DI({1'b0,Q[14:8]}),
        .O(D[15:8]),
        .S({\D16.DEL0[8].U_SRL_i_2__0_n_0 ,\D16.DEL0[8].U_SRL_i_3__0_n_0 ,\D16.DEL0[8].U_SRL_i_4__0_n_0 ,\D16.DEL0[8].U_SRL_i_5__0_n_0 ,\D16.DEL0[8].U_SRL_i_6__0_n_0 ,\D16.DEL0[8].U_SRL_i_7__0_n_0 ,\D16.DEL0[8].U_SRL_i_8__0_n_0 ,\D16.DEL0[8].U_SRL_i_9__0_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_2__0 
       (.I0(Q[15]),
        .I1(P[15]),
        .O(\D16.DEL0[8].U_SRL_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_3__0 
       (.I0(Q[14]),
        .I1(P[14]),
        .O(\D16.DEL0[8].U_SRL_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_4__0 
       (.I0(Q[13]),
        .I1(P[13]),
        .O(\D16.DEL0[8].U_SRL_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_5__0 
       (.I0(Q[12]),
        .I1(P[12]),
        .O(\D16.DEL0[8].U_SRL_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_6__0 
       (.I0(Q[11]),
        .I1(P[11]),
        .O(\D16.DEL0[8].U_SRL_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_7__0 
       (.I0(Q[10]),
        .I1(P[10]),
        .O(\D16.DEL0[8].U_SRL_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_8__0 
       (.I0(Q[9]),
        .I1(P[9]),
        .O(\D16.DEL0[8].U_SRL_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \D16.DEL0[8].U_SRL_i_9__0 
       (.I0(Q[8]),
        .I1(P[8]),
        .O(\D16.DEL0[8].U_SRL_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0 " *) 
  (* srl_name = "\activity_blocks[0].dutG/DZ2_78/D16.DEL0[9].U_SRL " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \D16.DEL0[9].U_SRL 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b1),
        .A3(1'b1),
        .CE(SE),
        .CLK(clk_i),
        .D(D[9]),
        .Q(clk_i_0[9]));
endmodule

(* ORIG_REF_NAME = "DualPortRAM" *) 
module switch_elements_DualPortRAM
   (ovDataOut_i,
    clk_i,
    rxd64_d3,
    \ovDataOut_reg[0] ,
    \ovDataOut_reg[63] ,
    \ovDataOut_reg[63]_0 ,
    \ovDataOut_reg[0]_0 );
  output [63:0]ovDataOut_i;
  input clk_i;
  input [63:0]rxd64_d3;
  input [6:0]\ovDataOut_reg[0] ;
  input [5:0]\ovDataOut_reg[63] ;
  input \ovDataOut_reg[63]_0 ;
  input \ovDataOut_reg[0]_0 ;

  wire clk_i;
  wire mem_reg_0_63_0_6_n_0;
  wire mem_reg_0_63_0_6_n_1;
  wire mem_reg_0_63_0_6_n_2;
  wire mem_reg_0_63_0_6_n_3;
  wire mem_reg_0_63_0_6_n_4;
  wire mem_reg_0_63_0_6_n_5;
  wire mem_reg_0_63_0_6_n_6;
  wire mem_reg_0_63_14_20_n_0;
  wire mem_reg_0_63_14_20_n_1;
  wire mem_reg_0_63_14_20_n_2;
  wire mem_reg_0_63_14_20_n_3;
  wire mem_reg_0_63_14_20_n_4;
  wire mem_reg_0_63_14_20_n_5;
  wire mem_reg_0_63_14_20_n_6;
  wire mem_reg_0_63_21_27_n_0;
  wire mem_reg_0_63_21_27_n_1;
  wire mem_reg_0_63_21_27_n_2;
  wire mem_reg_0_63_21_27_n_3;
  wire mem_reg_0_63_21_27_n_4;
  wire mem_reg_0_63_21_27_n_5;
  wire mem_reg_0_63_21_27_n_6;
  wire mem_reg_0_63_28_34_n_0;
  wire mem_reg_0_63_28_34_n_1;
  wire mem_reg_0_63_28_34_n_2;
  wire mem_reg_0_63_28_34_n_3;
  wire mem_reg_0_63_28_34_n_4;
  wire mem_reg_0_63_28_34_n_5;
  wire mem_reg_0_63_28_34_n_6;
  wire mem_reg_0_63_35_41_n_0;
  wire mem_reg_0_63_35_41_n_1;
  wire mem_reg_0_63_35_41_n_2;
  wire mem_reg_0_63_35_41_n_3;
  wire mem_reg_0_63_35_41_n_4;
  wire mem_reg_0_63_35_41_n_5;
  wire mem_reg_0_63_35_41_n_6;
  wire mem_reg_0_63_42_48_n_0;
  wire mem_reg_0_63_42_48_n_1;
  wire mem_reg_0_63_42_48_n_2;
  wire mem_reg_0_63_42_48_n_3;
  wire mem_reg_0_63_42_48_n_4;
  wire mem_reg_0_63_42_48_n_5;
  wire mem_reg_0_63_42_48_n_6;
  wire mem_reg_0_63_49_55_n_0;
  wire mem_reg_0_63_49_55_n_1;
  wire mem_reg_0_63_49_55_n_2;
  wire mem_reg_0_63_49_55_n_3;
  wire mem_reg_0_63_49_55_n_4;
  wire mem_reg_0_63_49_55_n_5;
  wire mem_reg_0_63_49_55_n_6;
  wire mem_reg_0_63_56_62_n_0;
  wire mem_reg_0_63_56_62_n_1;
  wire mem_reg_0_63_56_62_n_2;
  wire mem_reg_0_63_56_62_n_3;
  wire mem_reg_0_63_56_62_n_4;
  wire mem_reg_0_63_56_62_n_5;
  wire mem_reg_0_63_56_62_n_6;
  wire mem_reg_0_63_63_63_n_0;
  wire mem_reg_0_63_7_13_n_0;
  wire mem_reg_0_63_7_13_n_1;
  wire mem_reg_0_63_7_13_n_2;
  wire mem_reg_0_63_7_13_n_3;
  wire mem_reg_0_63_7_13_n_4;
  wire mem_reg_0_63_7_13_n_5;
  wire mem_reg_0_63_7_13_n_6;
  wire mem_reg_64_127_0_6_n_0;
  wire mem_reg_64_127_0_6_n_1;
  wire mem_reg_64_127_0_6_n_2;
  wire mem_reg_64_127_0_6_n_3;
  wire mem_reg_64_127_0_6_n_4;
  wire mem_reg_64_127_0_6_n_5;
  wire mem_reg_64_127_0_6_n_6;
  wire mem_reg_64_127_14_20_n_0;
  wire mem_reg_64_127_14_20_n_1;
  wire mem_reg_64_127_14_20_n_2;
  wire mem_reg_64_127_14_20_n_3;
  wire mem_reg_64_127_14_20_n_4;
  wire mem_reg_64_127_14_20_n_5;
  wire mem_reg_64_127_14_20_n_6;
  wire mem_reg_64_127_21_27_n_0;
  wire mem_reg_64_127_21_27_n_1;
  wire mem_reg_64_127_21_27_n_2;
  wire mem_reg_64_127_21_27_n_3;
  wire mem_reg_64_127_21_27_n_4;
  wire mem_reg_64_127_21_27_n_5;
  wire mem_reg_64_127_21_27_n_6;
  wire mem_reg_64_127_28_34_n_0;
  wire mem_reg_64_127_28_34_n_1;
  wire mem_reg_64_127_28_34_n_2;
  wire mem_reg_64_127_28_34_n_3;
  wire mem_reg_64_127_28_34_n_4;
  wire mem_reg_64_127_28_34_n_5;
  wire mem_reg_64_127_28_34_n_6;
  wire mem_reg_64_127_35_41_n_0;
  wire mem_reg_64_127_35_41_n_1;
  wire mem_reg_64_127_35_41_n_2;
  wire mem_reg_64_127_35_41_n_3;
  wire mem_reg_64_127_35_41_n_4;
  wire mem_reg_64_127_35_41_n_5;
  wire mem_reg_64_127_35_41_n_6;
  wire mem_reg_64_127_42_48_n_0;
  wire mem_reg_64_127_42_48_n_1;
  wire mem_reg_64_127_42_48_n_2;
  wire mem_reg_64_127_42_48_n_3;
  wire mem_reg_64_127_42_48_n_4;
  wire mem_reg_64_127_42_48_n_5;
  wire mem_reg_64_127_42_48_n_6;
  wire mem_reg_64_127_49_55_n_0;
  wire mem_reg_64_127_49_55_n_1;
  wire mem_reg_64_127_49_55_n_2;
  wire mem_reg_64_127_49_55_n_3;
  wire mem_reg_64_127_49_55_n_4;
  wire mem_reg_64_127_49_55_n_5;
  wire mem_reg_64_127_49_55_n_6;
  wire mem_reg_64_127_56_62_n_0;
  wire mem_reg_64_127_56_62_n_1;
  wire mem_reg_64_127_56_62_n_2;
  wire mem_reg_64_127_56_62_n_3;
  wire mem_reg_64_127_56_62_n_4;
  wire mem_reg_64_127_56_62_n_5;
  wire mem_reg_64_127_56_62_n_6;
  wire mem_reg_64_127_63_63_n_0;
  wire mem_reg_64_127_7_13_n_0;
  wire mem_reg_64_127_7_13_n_1;
  wire mem_reg_64_127_7_13_n_2;
  wire mem_reg_64_127_7_13_n_3;
  wire mem_reg_64_127_7_13_n_4;
  wire mem_reg_64_127_7_13_n_5;
  wire mem_reg_64_127_7_13_n_6;
  wire [63:0]ovDataOut_i;
  wire [6:0]\ovDataOut_reg[0] ;
  wire \ovDataOut_reg[0]_0 ;
  wire [5:0]\ovDataOut_reg[63] ;
  wire \ovDataOut_reg[63]_0 ;
  wire [63:0]rxd64_d3;
  wire NLW_mem_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_28_34_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_35_41_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_42_48_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_49_55_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_56_62_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_63_63_SPO_UNCONNECTED;
  wire NLW_mem_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_28_34_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_35_41_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_42_48_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_49_55_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_56_62_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_63_63_SPO_UNCONNECTED;
  wire NLW_mem_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD32714 mem_reg_0_63_0_6
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[0]),
        .DIB(rxd64_d3[1]),
        .DIC(rxd64_d3[2]),
        .DID(rxd64_d3[3]),
        .DIE(rxd64_d3[4]),
        .DIF(rxd64_d3[5]),
        .DIG(rxd64_d3[6]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_0_6_n_0),
        .DOB(mem_reg_0_63_0_6_n_1),
        .DOC(mem_reg_0_63_0_6_n_2),
        .DOD(mem_reg_0_63_0_6_n_3),
        .DOE(mem_reg_0_63_0_6_n_4),
        .DOF(mem_reg_0_63_0_6_n_5),
        .DOG(mem_reg_0_63_0_6_n_6),
        .DOH(NLW_mem_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD32715 mem_reg_0_63_14_20
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[14]),
        .DIB(rxd64_d3[15]),
        .DIC(rxd64_d3[16]),
        .DID(rxd64_d3[17]),
        .DIE(rxd64_d3[18]),
        .DIF(rxd64_d3[19]),
        .DIG(rxd64_d3[20]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_14_20_n_0),
        .DOB(mem_reg_0_63_14_20_n_1),
        .DOC(mem_reg_0_63_14_20_n_2),
        .DOD(mem_reg_0_63_14_20_n_3),
        .DOE(mem_reg_0_63_14_20_n_4),
        .DOF(mem_reg_0_63_14_20_n_5),
        .DOG(mem_reg_0_63_14_20_n_6),
        .DOH(NLW_mem_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD32716 mem_reg_0_63_21_27
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[21]),
        .DIB(rxd64_d3[22]),
        .DIC(rxd64_d3[23]),
        .DID(rxd64_d3[24]),
        .DIE(rxd64_d3[25]),
        .DIF(rxd64_d3[26]),
        .DIG(rxd64_d3[27]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_21_27_n_0),
        .DOB(mem_reg_0_63_21_27_n_1),
        .DOC(mem_reg_0_63_21_27_n_2),
        .DOD(mem_reg_0_63_21_27_n_3),
        .DOE(mem_reg_0_63_21_27_n_4),
        .DOF(mem_reg_0_63_21_27_n_5),
        .DOG(mem_reg_0_63_21_27_n_6),
        .DOH(NLW_mem_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "34" *) 
  RAM64M8_HD32717 mem_reg_0_63_28_34
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[28]),
        .DIB(rxd64_d3[29]),
        .DIC(rxd64_d3[30]),
        .DID(rxd64_d3[31]),
        .DIE(rxd64_d3[32]),
        .DIF(rxd64_d3[33]),
        .DIG(rxd64_d3[34]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_28_34_n_0),
        .DOB(mem_reg_0_63_28_34_n_1),
        .DOC(mem_reg_0_63_28_34_n_2),
        .DOD(mem_reg_0_63_28_34_n_3),
        .DOE(mem_reg_0_63_28_34_n_4),
        .DOF(mem_reg_0_63_28_34_n_5),
        .DOG(mem_reg_0_63_28_34_n_6),
        .DOH(NLW_mem_reg_0_63_28_34_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "35" *) 
  (* ram_slice_end = "41" *) 
  RAM64M8_HD32718 mem_reg_0_63_35_41
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[35]),
        .DIB(rxd64_d3[36]),
        .DIC(rxd64_d3[37]),
        .DID(rxd64_d3[38]),
        .DIE(rxd64_d3[39]),
        .DIF(rxd64_d3[40]),
        .DIG(rxd64_d3[41]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_35_41_n_0),
        .DOB(mem_reg_0_63_35_41_n_1),
        .DOC(mem_reg_0_63_35_41_n_2),
        .DOD(mem_reg_0_63_35_41_n_3),
        .DOE(mem_reg_0_63_35_41_n_4),
        .DOF(mem_reg_0_63_35_41_n_5),
        .DOG(mem_reg_0_63_35_41_n_6),
        .DOH(NLW_mem_reg_0_63_35_41_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "42" *) 
  (* ram_slice_end = "48" *) 
  RAM64M8_HD32719 mem_reg_0_63_42_48
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[42]),
        .DIB(rxd64_d3[43]),
        .DIC(rxd64_d3[44]),
        .DID(rxd64_d3[45]),
        .DIE(rxd64_d3[46]),
        .DIF(rxd64_d3[47]),
        .DIG(rxd64_d3[48]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_42_48_n_0),
        .DOB(mem_reg_0_63_42_48_n_1),
        .DOC(mem_reg_0_63_42_48_n_2),
        .DOD(mem_reg_0_63_42_48_n_3),
        .DOE(mem_reg_0_63_42_48_n_4),
        .DOF(mem_reg_0_63_42_48_n_5),
        .DOG(mem_reg_0_63_42_48_n_6),
        .DOH(NLW_mem_reg_0_63_42_48_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "49" *) 
  (* ram_slice_end = "55" *) 
  RAM64M8_HD32720 mem_reg_0_63_49_55
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[49]),
        .DIB(rxd64_d3[50]),
        .DIC(rxd64_d3[51]),
        .DID(rxd64_d3[52]),
        .DIE(rxd64_d3[53]),
        .DIF(rxd64_d3[54]),
        .DIG(rxd64_d3[55]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_49_55_n_0),
        .DOB(mem_reg_0_63_49_55_n_1),
        .DOC(mem_reg_0_63_49_55_n_2),
        .DOD(mem_reg_0_63_49_55_n_3),
        .DOE(mem_reg_0_63_49_55_n_4),
        .DOF(mem_reg_0_63_49_55_n_5),
        .DOG(mem_reg_0_63_49_55_n_6),
        .DOH(NLW_mem_reg_0_63_49_55_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "56" *) 
  (* ram_slice_end = "62" *) 
  RAM64M8_HD32721 mem_reg_0_63_56_62
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[56]),
        .DIB(rxd64_d3[57]),
        .DIC(rxd64_d3[58]),
        .DID(rxd64_d3[59]),
        .DIE(rxd64_d3[60]),
        .DIF(rxd64_d3[61]),
        .DIG(rxd64_d3[62]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_56_62_n_0),
        .DOB(mem_reg_0_63_56_62_n_1),
        .DOC(mem_reg_0_63_56_62_n_2),
        .DOD(mem_reg_0_63_56_62_n_3),
        .DOE(mem_reg_0_63_56_62_n_4),
        .DOF(mem_reg_0_63_56_62_n_5),
        .DOG(mem_reg_0_63_56_62_n_6),
        .DOH(NLW_mem_reg_0_63_56_62_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT = "64'h0000000000000000" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "63" *) 
  (* ram_slice_end = "63" *) 
  RAM64X1D_HD32722 mem_reg_0_63_63_63
       (.A0(\ovDataOut_reg[63] [0]),
        .A1(\ovDataOut_reg[63] [1]),
        .A2(\ovDataOut_reg[63] [2]),
        .A3(\ovDataOut_reg[63] [3]),
        .A4(\ovDataOut_reg[63] [4]),
        .A5(\ovDataOut_reg[63] [5]),
        .D(rxd64_d3[63]),
        .DPO(mem_reg_0_63_63_63_n_0),
        .DPRA0(\ovDataOut_reg[0] [0]),
        .DPRA1(\ovDataOut_reg[0] [1]),
        .DPRA2(\ovDataOut_reg[0] [2]),
        .DPRA3(\ovDataOut_reg[0] [3]),
        .DPRA4(\ovDataOut_reg[0] [4]),
        .DPRA5(\ovDataOut_reg[0] [5]),
        .SPO(NLW_mem_reg_0_63_63_63_SPO_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD32723 mem_reg_0_63_7_13
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[7]),
        .DIB(rxd64_d3[8]),
        .DIC(rxd64_d3[9]),
        .DID(rxd64_d3[10]),
        .DIE(rxd64_d3[11]),
        .DIF(rxd64_d3[12]),
        .DIG(rxd64_d3[13]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_7_13_n_0),
        .DOB(mem_reg_0_63_7_13_n_1),
        .DOC(mem_reg_0_63_7_13_n_2),
        .DOD(mem_reg_0_63_7_13_n_3),
        .DOE(mem_reg_0_63_7_13_n_4),
        .DOF(mem_reg_0_63_7_13_n_5),
        .DOG(mem_reg_0_63_7_13_n_6),
        .DOH(NLW_mem_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[63]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD32724 mem_reg_64_127_0_6
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[0]),
        .DIB(rxd64_d3[1]),
        .DIC(rxd64_d3[2]),
        .DID(rxd64_d3[3]),
        .DIE(rxd64_d3[4]),
        .DIF(rxd64_d3[5]),
        .DIG(rxd64_d3[6]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_0_6_n_0),
        .DOB(mem_reg_64_127_0_6_n_1),
        .DOC(mem_reg_64_127_0_6_n_2),
        .DOD(mem_reg_64_127_0_6_n_3),
        .DOE(mem_reg_64_127_0_6_n_4),
        .DOF(mem_reg_64_127_0_6_n_5),
        .DOG(mem_reg_64_127_0_6_n_6),
        .DOH(NLW_mem_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD32725 mem_reg_64_127_14_20
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[14]),
        .DIB(rxd64_d3[15]),
        .DIC(rxd64_d3[16]),
        .DID(rxd64_d3[17]),
        .DIE(rxd64_d3[18]),
        .DIF(rxd64_d3[19]),
        .DIG(rxd64_d3[20]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_14_20_n_0),
        .DOB(mem_reg_64_127_14_20_n_1),
        .DOC(mem_reg_64_127_14_20_n_2),
        .DOD(mem_reg_64_127_14_20_n_3),
        .DOE(mem_reg_64_127_14_20_n_4),
        .DOF(mem_reg_64_127_14_20_n_5),
        .DOG(mem_reg_64_127_14_20_n_6),
        .DOH(NLW_mem_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD32726 mem_reg_64_127_21_27
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[21]),
        .DIB(rxd64_d3[22]),
        .DIC(rxd64_d3[23]),
        .DID(rxd64_d3[24]),
        .DIE(rxd64_d3[25]),
        .DIF(rxd64_d3[26]),
        .DIG(rxd64_d3[27]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_21_27_n_0),
        .DOB(mem_reg_64_127_21_27_n_1),
        .DOC(mem_reg_64_127_21_27_n_2),
        .DOD(mem_reg_64_127_21_27_n_3),
        .DOE(mem_reg_64_127_21_27_n_4),
        .DOF(mem_reg_64_127_21_27_n_5),
        .DOG(mem_reg_64_127_21_27_n_6),
        .DOH(NLW_mem_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "34" *) 
  RAM64M8_HD32727 mem_reg_64_127_28_34
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[28]),
        .DIB(rxd64_d3[29]),
        .DIC(rxd64_d3[30]),
        .DID(rxd64_d3[31]),
        .DIE(rxd64_d3[32]),
        .DIF(rxd64_d3[33]),
        .DIG(rxd64_d3[34]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_28_34_n_0),
        .DOB(mem_reg_64_127_28_34_n_1),
        .DOC(mem_reg_64_127_28_34_n_2),
        .DOD(mem_reg_64_127_28_34_n_3),
        .DOE(mem_reg_64_127_28_34_n_4),
        .DOF(mem_reg_64_127_28_34_n_5),
        .DOG(mem_reg_64_127_28_34_n_6),
        .DOH(NLW_mem_reg_64_127_28_34_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "35" *) 
  (* ram_slice_end = "41" *) 
  RAM64M8_HD32728 mem_reg_64_127_35_41
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[35]),
        .DIB(rxd64_d3[36]),
        .DIC(rxd64_d3[37]),
        .DID(rxd64_d3[38]),
        .DIE(rxd64_d3[39]),
        .DIF(rxd64_d3[40]),
        .DIG(rxd64_d3[41]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_35_41_n_0),
        .DOB(mem_reg_64_127_35_41_n_1),
        .DOC(mem_reg_64_127_35_41_n_2),
        .DOD(mem_reg_64_127_35_41_n_3),
        .DOE(mem_reg_64_127_35_41_n_4),
        .DOF(mem_reg_64_127_35_41_n_5),
        .DOG(mem_reg_64_127_35_41_n_6),
        .DOH(NLW_mem_reg_64_127_35_41_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "42" *) 
  (* ram_slice_end = "48" *) 
  RAM64M8_HD32729 mem_reg_64_127_42_48
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[42]),
        .DIB(rxd64_d3[43]),
        .DIC(rxd64_d3[44]),
        .DID(rxd64_d3[45]),
        .DIE(rxd64_d3[46]),
        .DIF(rxd64_d3[47]),
        .DIG(rxd64_d3[48]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_42_48_n_0),
        .DOB(mem_reg_64_127_42_48_n_1),
        .DOC(mem_reg_64_127_42_48_n_2),
        .DOD(mem_reg_64_127_42_48_n_3),
        .DOE(mem_reg_64_127_42_48_n_4),
        .DOF(mem_reg_64_127_42_48_n_5),
        .DOG(mem_reg_64_127_42_48_n_6),
        .DOH(NLW_mem_reg_64_127_42_48_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "49" *) 
  (* ram_slice_end = "55" *) 
  RAM64M8_HD32730 mem_reg_64_127_49_55
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[49]),
        .DIB(rxd64_d3[50]),
        .DIC(rxd64_d3[51]),
        .DID(rxd64_d3[52]),
        .DIE(rxd64_d3[53]),
        .DIF(rxd64_d3[54]),
        .DIG(rxd64_d3[55]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_49_55_n_0),
        .DOB(mem_reg_64_127_49_55_n_1),
        .DOC(mem_reg_64_127_49_55_n_2),
        .DOD(mem_reg_64_127_49_55_n_3),
        .DOE(mem_reg_64_127_49_55_n_4),
        .DOF(mem_reg_64_127_49_55_n_5),
        .DOG(mem_reg_64_127_49_55_n_6),
        .DOH(NLW_mem_reg_64_127_49_55_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "56" *) 
  (* ram_slice_end = "62" *) 
  RAM64M8_HD32731 mem_reg_64_127_56_62
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[56]),
        .DIB(rxd64_d3[57]),
        .DIC(rxd64_d3[58]),
        .DID(rxd64_d3[59]),
        .DIE(rxd64_d3[60]),
        .DIF(rxd64_d3[61]),
        .DIG(rxd64_d3[62]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_56_62_n_0),
        .DOB(mem_reg_64_127_56_62_n_1),
        .DOC(mem_reg_64_127_56_62_n_2),
        .DOD(mem_reg_64_127_56_62_n_3),
        .DOE(mem_reg_64_127_56_62_n_4),
        .DOF(mem_reg_64_127_56_62_n_5),
        .DOG(mem_reg_64_127_56_62_n_6),
        .DOH(NLW_mem_reg_64_127_56_62_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT = "64'h0000000000000000" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "63" *) 
  (* ram_slice_end = "63" *) 
  RAM64X1D_HD32732 mem_reg_64_127_63_63
       (.A0(\ovDataOut_reg[63] [0]),
        .A1(\ovDataOut_reg[63] [1]),
        .A2(\ovDataOut_reg[63] [2]),
        .A3(\ovDataOut_reg[63] [3]),
        .A4(\ovDataOut_reg[63] [4]),
        .A5(\ovDataOut_reg[63] [5]),
        .D(rxd64_d3[63]),
        .DPO(mem_reg_64_127_63_63_n_0),
        .DPRA0(\ovDataOut_reg[0] [0]),
        .DPRA1(\ovDataOut_reg[0] [1]),
        .DPRA2(\ovDataOut_reg[0] [2]),
        .DPRA3(\ovDataOut_reg[0] [3]),
        .DPRA4(\ovDataOut_reg[0] [4]),
        .DPRA5(\ovDataOut_reg[0] [5]),
        .SPO(NLW_mem_reg_64_127_63_63_SPO_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "8192" *) 
  (* RTL_RAM_NAME = "datapath_main/rxdatain/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD32733 mem_reg_64_127_7_13
       (.ADDRA(\ovDataOut_reg[0] [5:0]),
        .ADDRB(\ovDataOut_reg[0] [5:0]),
        .ADDRC(\ovDataOut_reg[0] [5:0]),
        .ADDRD(\ovDataOut_reg[0] [5:0]),
        .ADDRE(\ovDataOut_reg[0] [5:0]),
        .ADDRF(\ovDataOut_reg[0] [5:0]),
        .ADDRG(\ovDataOut_reg[0] [5:0]),
        .ADDRH(\ovDataOut_reg[63] ),
        .DIA(rxd64_d3[7]),
        .DIB(rxd64_d3[8]),
        .DIC(rxd64_d3[9]),
        .DID(rxd64_d3[10]),
        .DIE(rxd64_d3[11]),
        .DIF(rxd64_d3[12]),
        .DIG(rxd64_d3[13]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_7_13_n_0),
        .DOB(mem_reg_64_127_7_13_n_1),
        .DOC(mem_reg_64_127_7_13_n_2),
        .DOD(mem_reg_64_127_7_13_n_3),
        .DOE(mem_reg_64_127_7_13_n_4),
        .DOF(mem_reg_64_127_7_13_n_5),
        .DOG(mem_reg_64_127_7_13_n_6),
        .DOH(NLW_mem_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[0]_i_1 
       (.I0(mem_reg_64_127_0_6_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_0),
        .O(ovDataOut_i[0]));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[10]_i_1 
       (.I0(mem_reg_64_127_7_13_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_3),
        .O(ovDataOut_i[10]));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[11]_i_1 
       (.I0(mem_reg_64_127_7_13_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_4),
        .O(ovDataOut_i[11]));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[12]_i_1 
       (.I0(mem_reg_64_127_7_13_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_5),
        .O(ovDataOut_i[12]));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[13]_i_1 
       (.I0(mem_reg_64_127_7_13_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_6),
        .O(ovDataOut_i[13]));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[14]_i_1 
       (.I0(mem_reg_64_127_14_20_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_0),
        .O(ovDataOut_i[14]));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[15]_i_1 
       (.I0(mem_reg_64_127_14_20_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_1),
        .O(ovDataOut_i[15]));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[16]_i_1 
       (.I0(mem_reg_64_127_14_20_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_2),
        .O(ovDataOut_i[16]));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[17]_i_1 
       (.I0(mem_reg_64_127_14_20_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_3),
        .O(ovDataOut_i[17]));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[18]_i_1 
       (.I0(mem_reg_64_127_14_20_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_4),
        .O(ovDataOut_i[18]));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[19]_i_1 
       (.I0(mem_reg_64_127_14_20_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_5),
        .O(ovDataOut_i[19]));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[1]_i_1 
       (.I0(mem_reg_64_127_0_6_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_1),
        .O(ovDataOut_i[1]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[20]_i_1 
       (.I0(mem_reg_64_127_14_20_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_14_20_n_6),
        .O(ovDataOut_i[20]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[21]_i_1 
       (.I0(mem_reg_64_127_21_27_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_0),
        .O(ovDataOut_i[21]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[22]_i_1 
       (.I0(mem_reg_64_127_21_27_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_1),
        .O(ovDataOut_i[22]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[23]_i_1 
       (.I0(mem_reg_64_127_21_27_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_2),
        .O(ovDataOut_i[23]));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[24]_i_1 
       (.I0(mem_reg_64_127_21_27_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_3),
        .O(ovDataOut_i[24]));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[25]_i_1 
       (.I0(mem_reg_64_127_21_27_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_4),
        .O(ovDataOut_i[25]));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[26]_i_1 
       (.I0(mem_reg_64_127_21_27_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_5),
        .O(ovDataOut_i[26]));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[27]_i_1 
       (.I0(mem_reg_64_127_21_27_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_21_27_n_6),
        .O(ovDataOut_i[27]));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[28]_i_1 
       (.I0(mem_reg_64_127_28_34_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_0),
        .O(ovDataOut_i[28]));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[29]_i_1 
       (.I0(mem_reg_64_127_28_34_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_1),
        .O(ovDataOut_i[29]));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[2]_i_1 
       (.I0(mem_reg_64_127_0_6_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_2),
        .O(ovDataOut_i[2]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[30]_i_1 
       (.I0(mem_reg_64_127_28_34_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_2),
        .O(ovDataOut_i[30]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[31]_i_1 
       (.I0(mem_reg_64_127_28_34_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_3),
        .O(ovDataOut_i[31]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[32]_i_1 
       (.I0(mem_reg_64_127_28_34_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_4),
        .O(ovDataOut_i[32]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[33]_i_1 
       (.I0(mem_reg_64_127_28_34_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_5),
        .O(ovDataOut_i[33]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[34]_i_1 
       (.I0(mem_reg_64_127_28_34_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_28_34_n_6),
        .O(ovDataOut_i[34]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[35]_i_1 
       (.I0(mem_reg_64_127_35_41_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_0),
        .O(ovDataOut_i[35]));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[36]_i_1 
       (.I0(mem_reg_64_127_35_41_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_1),
        .O(ovDataOut_i[36]));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[37]_i_1 
       (.I0(mem_reg_64_127_35_41_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_2),
        .O(ovDataOut_i[37]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[38]_i_1 
       (.I0(mem_reg_64_127_35_41_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_3),
        .O(ovDataOut_i[38]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[39]_i_1 
       (.I0(mem_reg_64_127_35_41_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_4),
        .O(ovDataOut_i[39]));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[3]_i_1 
       (.I0(mem_reg_64_127_0_6_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_3),
        .O(ovDataOut_i[3]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[40]_i_1 
       (.I0(mem_reg_64_127_35_41_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_5),
        .O(ovDataOut_i[40]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[41]_i_1 
       (.I0(mem_reg_64_127_35_41_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_35_41_n_6),
        .O(ovDataOut_i[41]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[42]_i_1 
       (.I0(mem_reg_64_127_42_48_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_0),
        .O(ovDataOut_i[42]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[43]_i_1 
       (.I0(mem_reg_64_127_42_48_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_1),
        .O(ovDataOut_i[43]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[44]_i_1 
       (.I0(mem_reg_64_127_42_48_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_2),
        .O(ovDataOut_i[44]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[45]_i_1 
       (.I0(mem_reg_64_127_42_48_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_3),
        .O(ovDataOut_i[45]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[46]_i_1 
       (.I0(mem_reg_64_127_42_48_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_4),
        .O(ovDataOut_i[46]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[47]_i_1 
       (.I0(mem_reg_64_127_42_48_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_5),
        .O(ovDataOut_i[47]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[48]_i_1 
       (.I0(mem_reg_64_127_42_48_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_42_48_n_6),
        .O(ovDataOut_i[48]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[49]_i_1 
       (.I0(mem_reg_64_127_49_55_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_0),
        .O(ovDataOut_i[49]));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[4]_i_1 
       (.I0(mem_reg_64_127_0_6_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_4),
        .O(ovDataOut_i[4]));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[50]_i_1 
       (.I0(mem_reg_64_127_49_55_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_1),
        .O(ovDataOut_i[50]));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[51]_i_1 
       (.I0(mem_reg_64_127_49_55_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_2),
        .O(ovDataOut_i[51]));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[52]_i_1 
       (.I0(mem_reg_64_127_49_55_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_3),
        .O(ovDataOut_i[52]));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[53]_i_1 
       (.I0(mem_reg_64_127_49_55_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_4),
        .O(ovDataOut_i[53]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[54]_i_1 
       (.I0(mem_reg_64_127_49_55_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_5),
        .O(ovDataOut_i[54]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[55]_i_1 
       (.I0(mem_reg_64_127_49_55_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_49_55_n_6),
        .O(ovDataOut_i[55]));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[56]_i_1 
       (.I0(mem_reg_64_127_56_62_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_0),
        .O(ovDataOut_i[56]));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[57]_i_1 
       (.I0(mem_reg_64_127_56_62_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_1),
        .O(ovDataOut_i[57]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[58]_i_1 
       (.I0(mem_reg_64_127_56_62_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_2),
        .O(ovDataOut_i[58]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[59]_i_1 
       (.I0(mem_reg_64_127_56_62_n_3),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_3),
        .O(ovDataOut_i[59]));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[5]_i_1 
       (.I0(mem_reg_64_127_0_6_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_5),
        .O(ovDataOut_i[5]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[60]_i_1 
       (.I0(mem_reg_64_127_56_62_n_4),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_4),
        .O(ovDataOut_i[60]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[61]_i_1 
       (.I0(mem_reg_64_127_56_62_n_5),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_5),
        .O(ovDataOut_i[61]));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[62]_i_1 
       (.I0(mem_reg_64_127_56_62_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_56_62_n_6),
        .O(ovDataOut_i[62]));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[63]_i_2 
       (.I0(mem_reg_64_127_63_63_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_63_63_n_0),
        .O(ovDataOut_i[63]));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[6]_i_1 
       (.I0(mem_reg_64_127_0_6_n_6),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_0_6_n_6),
        .O(ovDataOut_i[6]));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[7]_i_1 
       (.I0(mem_reg_64_127_7_13_n_0),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_0),
        .O(ovDataOut_i[7]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[8]_i_1 
       (.I0(mem_reg_64_127_7_13_n_1),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_1),
        .O(ovDataOut_i[8]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[9]_i_1 
       (.I0(mem_reg_64_127_7_13_n_2),
        .I1(\ovDataOut_reg[0] [6]),
        .I2(mem_reg_0_63_7_13_n_2),
        .O(ovDataOut_i[9]));
endmodule

(* ORIG_REF_NAME = "DualPortRAM_ASYN" *) 
module switch_elements_DualPortRAM_ASYN
   (clk_i_0,
    clk_i,
    E,
    MemDataIn,
    ADDRH,
    D);
  output [71:0]clk_i_0;
  input clk_i;
  input [0:0]E;
  input [71:0]MemDataIn;
  input [4:0]ADDRH;
  input [4:0]D;

  wire [4:0]ADDRH;
  wire [4:0]D;
  wire [0:0]E;
  wire [71:0]MemDataIn;
  wire clk_i;
  wire [71:0]clk_i_0;
  wire \qvRAddr_reg_n_0_[0] ;
  wire \qvRAddr_reg_n_0_[1] ;
  wire \qvRAddr_reg_n_0_[2] ;
  wire \qvRAddr_reg_n_0_[3] ;
  wire \qvRAddr_reg_n_0_[4] ;
  wire [1:0]NLW_mem_reg_0_31_0_13_DOH_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_14_27_DOH_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_28_41_DOH_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_42_55_DOH_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_56_69_DOH_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOB_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOC_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOD_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOE_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOF_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOG_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_31_70_71_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "2304" *) 
  (* RTL_RAM_NAME = "rx_rs/datapath/RealignInst/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "31" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "13" *) 
  RAM32M16_HD32734 mem_reg_0_31_0_13
       (.ADDRA({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRB({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRC({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRD({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRE({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRF({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRG({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRH(ADDRH),
        .DIA(MemDataIn[1:0]),
        .DIB(MemDataIn[3:2]),
        .DIC(MemDataIn[5:4]),
        .DID(MemDataIn[7:6]),
        .DIE(MemDataIn[9:8]),
        .DIF(MemDataIn[11:10]),
        .DIG(MemDataIn[13:12]),
        .DIH({1'b0,1'b0}),
        .DOA(clk_i_0[1:0]),
        .DOB(clk_i_0[3:2]),
        .DOC(clk_i_0[5:4]),
        .DOD(clk_i_0[7:6]),
        .DOE(clk_i_0[9:8]),
        .DOF(clk_i_0[11:10]),
        .DOG(clk_i_0[13:12]),
        .DOH(NLW_mem_reg_0_31_0_13_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(E));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "2304" *) 
  (* RTL_RAM_NAME = "rx_rs/datapath/RealignInst/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "31" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "27" *) 
  RAM32M16_HD32735 mem_reg_0_31_14_27
       (.ADDRA({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRB({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRC({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRD({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRE({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRF({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRG({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRH(ADDRH),
        .DIA(MemDataIn[15:14]),
        .DIB(MemDataIn[17:16]),
        .DIC(MemDataIn[19:18]),
        .DID(MemDataIn[21:20]),
        .DIE(MemDataIn[23:22]),
        .DIF(MemDataIn[25:24]),
        .DIG(MemDataIn[27:26]),
        .DIH({1'b0,1'b0}),
        .DOA(clk_i_0[15:14]),
        .DOB(clk_i_0[17:16]),
        .DOC(clk_i_0[19:18]),
        .DOD(clk_i_0[21:20]),
        .DOE(clk_i_0[23:22]),
        .DOF(clk_i_0[25:24]),
        .DOG(clk_i_0[27:26]),
        .DOH(NLW_mem_reg_0_31_14_27_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(E));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "2304" *) 
  (* RTL_RAM_NAME = "rx_rs/datapath/RealignInst/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "31" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "41" *) 
  RAM32M16_HD32736 mem_reg_0_31_28_41
       (.ADDRA({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRB({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRC({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRD({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRE({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRF({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRG({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRH(ADDRH),
        .DIA(MemDataIn[29:28]),
        .DIB(MemDataIn[31:30]),
        .DIC(MemDataIn[33:32]),
        .DID(MemDataIn[35:34]),
        .DIE(MemDataIn[37:36]),
        .DIF(MemDataIn[39:38]),
        .DIG(MemDataIn[41:40]),
        .DIH({1'b0,1'b0}),
        .DOA(clk_i_0[29:28]),
        .DOB(clk_i_0[31:30]),
        .DOC(clk_i_0[33:32]),
        .DOD(clk_i_0[35:34]),
        .DOE(clk_i_0[37:36]),
        .DOF(clk_i_0[39:38]),
        .DOG(clk_i_0[41:40]),
        .DOH(NLW_mem_reg_0_31_28_41_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(E));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "2304" *) 
  (* RTL_RAM_NAME = "rx_rs/datapath/RealignInst/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "31" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "42" *) 
  (* ram_slice_end = "55" *) 
  RAM32M16_HD32737 mem_reg_0_31_42_55
       (.ADDRA({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRB({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRC({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRD({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRE({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRF({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRG({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRH(ADDRH),
        .DIA(MemDataIn[43:42]),
        .DIB(MemDataIn[45:44]),
        .DIC(MemDataIn[47:46]),
        .DID(MemDataIn[49:48]),
        .DIE(MemDataIn[51:50]),
        .DIF(MemDataIn[53:52]),
        .DIG(MemDataIn[55:54]),
        .DIH({1'b0,1'b0}),
        .DOA(clk_i_0[43:42]),
        .DOB(clk_i_0[45:44]),
        .DOC(clk_i_0[47:46]),
        .DOD(clk_i_0[49:48]),
        .DOE(clk_i_0[51:50]),
        .DOF(clk_i_0[53:52]),
        .DOG(clk_i_0[55:54]),
        .DOH(NLW_mem_reg_0_31_42_55_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(E));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "2304" *) 
  (* RTL_RAM_NAME = "rx_rs/datapath/RealignInst/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "31" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "56" *) 
  (* ram_slice_end = "69" *) 
  RAM32M16_HD32738 mem_reg_0_31_56_69
       (.ADDRA({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRB({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRC({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRD({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRE({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRF({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRG({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRH(ADDRH),
        .DIA(MemDataIn[57:56]),
        .DIB(MemDataIn[59:58]),
        .DIC(MemDataIn[61:60]),
        .DID(MemDataIn[63:62]),
        .DIE(MemDataIn[65:64]),
        .DIF(MemDataIn[67:66]),
        .DIG(MemDataIn[69:68]),
        .DIH({1'b0,1'b0}),
        .DOA(clk_i_0[57:56]),
        .DOB(clk_i_0[59:58]),
        .DOC(clk_i_0[61:60]),
        .DOD(clk_i_0[63:62]),
        .DOE(clk_i_0[65:64]),
        .DOF(clk_i_0[67:66]),
        .DOG(clk_i_0[69:68]),
        .DOH(NLW_mem_reg_0_31_56_69_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(E));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "2304" *) 
  (* RTL_RAM_NAME = "rx_rs/datapath/RealignInst/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "31" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "70" *) 
  (* ram_slice_end = "71" *) 
  RAM32M16_HD32739 mem_reg_0_31_70_71
       (.ADDRA({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRB({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRC({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRD({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRE({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRF({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRG({\qvRAddr_reg_n_0_[4] ,\qvRAddr_reg_n_0_[3] ,\qvRAddr_reg_n_0_[2] ,\qvRAddr_reg_n_0_[1] ,\qvRAddr_reg_n_0_[0] }),
        .ADDRH(ADDRH),
        .DIA(MemDataIn[71:70]),
        .DIB({1'b0,1'b0}),
        .DIC({1'b0,1'b0}),
        .DID({1'b0,1'b0}),
        .DIE({1'b0,1'b0}),
        .DIF({1'b0,1'b0}),
        .DIG({1'b0,1'b0}),
        .DIH({1'b0,1'b0}),
        .DOA(clk_i_0[71:70]),
        .DOB(NLW_mem_reg_0_31_70_71_DOB_UNCONNECTED[1:0]),
        .DOC(NLW_mem_reg_0_31_70_71_DOC_UNCONNECTED[1:0]),
        .DOD(NLW_mem_reg_0_31_70_71_DOD_UNCONNECTED[1:0]),
        .DOE(NLW_mem_reg_0_31_70_71_DOE_UNCONNECTED[1:0]),
        .DOF(NLW_mem_reg_0_31_70_71_DOF_UNCONNECTED[1:0]),
        .DOG(NLW_mem_reg_0_31_70_71_DOG_UNCONNECTED[1:0]),
        .DOH(NLW_mem_reg_0_31_70_71_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(E));
  FDRE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(D[0]),
        .Q(\qvRAddr_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(D[1]),
        .Q(\qvRAddr_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(D[2]),
        .Q(\qvRAddr_reg_n_0_[2] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(D[3]),
        .Q(\qvRAddr_reg_n_0_[3] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(D[4]),
        .Q(\qvRAddr_reg_n_0_[4] ),
        .R(1'b0));
endmodule

(* ORIG_REF_NAME = "DualPortRAM" *) 
module switch_elements_DualPortRAM__parameterized0
   (ovDataOut_i,
    clk_i,
    vDataIn,
    Q,
    \ovDataOut_reg[7] ,
    \ovDataOut_reg[0] ,
    \ovDataOut_reg[7]_0 );
  output [7:0]ovDataOut_i;
  input clk_i;
  input [7:0]vDataIn;
  input [6:0]Q;
  input [5:0]\ovDataOut_reg[7] ;
  input \ovDataOut_reg[0] ;
  input \ovDataOut_reg[7]_0 ;

  wire [6:0]Q;
  wire clk_i;
  wire mem_reg_0_63_0_6_n_0;
  wire mem_reg_0_63_0_6_n_1;
  wire mem_reg_0_63_0_6_n_2;
  wire mem_reg_0_63_0_6_n_3;
  wire mem_reg_0_63_0_6_n_4;
  wire mem_reg_0_63_0_6_n_5;
  wire mem_reg_0_63_0_6_n_6;
  wire mem_reg_0_63_7_7_n_0;
  wire mem_reg_64_127_0_6_n_0;
  wire mem_reg_64_127_0_6_n_1;
  wire mem_reg_64_127_0_6_n_2;
  wire mem_reg_64_127_0_6_n_3;
  wire mem_reg_64_127_0_6_n_4;
  wire mem_reg_64_127_0_6_n_5;
  wire mem_reg_64_127_0_6_n_6;
  wire mem_reg_64_127_7_7_n_0;
  wire [7:0]ovDataOut_i;
  wire \ovDataOut_reg[0] ;
  wire [5:0]\ovDataOut_reg[7] ;
  wire \ovDataOut_reg[7]_0 ;
  wire [7:0]vDataIn;
  wire NLW_mem_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_mem_reg_0_63_7_7_SPO_UNCONNECTED;
  wire NLW_mem_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_mem_reg_64_127_7_7_SPO_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "1024" *) 
  (* RTL_RAM_NAME = "datapath_main/rxcntrlin/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_UNIQ_BASE_ mem_reg_0_63_0_6
       (.ADDRA(Q[5:0]),
        .ADDRB(Q[5:0]),
        .ADDRC(Q[5:0]),
        .ADDRD(Q[5:0]),
        .ADDRE(Q[5:0]),
        .ADDRF(Q[5:0]),
        .ADDRG(Q[5:0]),
        .ADDRH(\ovDataOut_reg[7] ),
        .DIA(vDataIn[0]),
        .DIB(vDataIn[1]),
        .DIC(vDataIn[2]),
        .DID(vDataIn[3]),
        .DIE(vDataIn[4]),
        .DIF(vDataIn[5]),
        .DIG(vDataIn[6]),
        .DIH(1'b0),
        .DOA(mem_reg_0_63_0_6_n_0),
        .DOB(mem_reg_0_63_0_6_n_1),
        .DOC(mem_reg_0_63_0_6_n_2),
        .DOD(mem_reg_0_63_0_6_n_3),
        .DOE(mem_reg_0_63_0_6_n_4),
        .DOF(mem_reg_0_63_0_6_n_5),
        .DOG(mem_reg_0_63_0_6_n_6),
        .DOH(NLW_mem_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0] ));
  (* INIT = "64'h0000000000000000" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "7" *) 
  RAM64X1D_UNIQ_BASE_ mem_reg_0_63_7_7
       (.A0(\ovDataOut_reg[7] [0]),
        .A1(\ovDataOut_reg[7] [1]),
        .A2(\ovDataOut_reg[7] [2]),
        .A3(\ovDataOut_reg[7] [3]),
        .A4(\ovDataOut_reg[7] [4]),
        .A5(\ovDataOut_reg[7] [5]),
        .D(vDataIn[7]),
        .DPO(mem_reg_0_63_7_7_n_0),
        .DPRA0(Q[0]),
        .DPRA1(Q[1]),
        .DPRA2(Q[2]),
        .DPRA3(Q[3]),
        .DPRA4(Q[4]),
        .DPRA5(Q[5]),
        .SPO(NLW_mem_reg_0_63_7_7_SPO_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[0] ));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "1024" *) 
  (* RTL_RAM_NAME = "datapath_main/rxcntrlin/Fifo_Storage/mem" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD32712 mem_reg_64_127_0_6
       (.ADDRA(Q[5:0]),
        .ADDRB(Q[5:0]),
        .ADDRC(Q[5:0]),
        .ADDRD(Q[5:0]),
        .ADDRE(Q[5:0]),
        .ADDRF(Q[5:0]),
        .ADDRG(Q[5:0]),
        .ADDRH(\ovDataOut_reg[7] ),
        .DIA(vDataIn[0]),
        .DIB(vDataIn[1]),
        .DIC(vDataIn[2]),
        .DID(vDataIn[3]),
        .DIE(vDataIn[4]),
        .DIF(vDataIn[5]),
        .DIG(vDataIn[6]),
        .DIH(1'b0),
        .DOA(mem_reg_64_127_0_6_n_0),
        .DOB(mem_reg_64_127_0_6_n_1),
        .DOC(mem_reg_64_127_0_6_n_2),
        .DOD(mem_reg_64_127_0_6_n_3),
        .DOE(mem_reg_64_127_0_6_n_4),
        .DOF(mem_reg_64_127_0_6_n_5),
        .DOG(mem_reg_64_127_0_6_n_6),
        .DOH(NLW_mem_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[7]_0 ));
  (* INIT = "64'h0000000000000000" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "7" *) 
  RAM64X1D_HD32713 mem_reg_64_127_7_7
       (.A0(\ovDataOut_reg[7] [0]),
        .A1(\ovDataOut_reg[7] [1]),
        .A2(\ovDataOut_reg[7] [2]),
        .A3(\ovDataOut_reg[7] [3]),
        .A4(\ovDataOut_reg[7] [4]),
        .A5(\ovDataOut_reg[7] [5]),
        .D(vDataIn[7]),
        .DPO(mem_reg_64_127_7_7_n_0),
        .DPRA0(Q[0]),
        .DPRA1(Q[1]),
        .DPRA2(Q[2]),
        .DPRA3(Q[3]),
        .DPRA4(Q[4]),
        .DPRA5(Q[5]),
        .SPO(NLW_mem_reg_64_127_7_7_SPO_UNCONNECTED),
        .WCLK(clk_i),
        .WE(\ovDataOut_reg[7]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[0]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_0),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_0),
        .O(ovDataOut_i[0]));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[1]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_1),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_1),
        .O(ovDataOut_i[1]));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[2]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_2),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_2),
        .O(ovDataOut_i[2]));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[3]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_3),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_3),
        .O(ovDataOut_i[3]));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[4]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_4),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_4),
        .O(ovDataOut_i[4]));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[5]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_5),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_5),
        .O(ovDataOut_i[5]));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[6]_i_1__0 
       (.I0(mem_reg_64_127_0_6_n_6),
        .I1(Q[6]),
        .I2(mem_reg_0_63_0_6_n_6),
        .O(ovDataOut_i[6]));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ovDataOut[7]_i_2 
       (.I0(mem_reg_64_127_7_7_n_0),
        .I1(Q[6]),
        .I2(mem_reg_0_63_7_7_n_0),
        .O(ovDataOut_i[7]));
endmodule

(* ORIG_REF_NAME = "FifoControl" *) 
module switch_elements_FifoControl
   (qEmpty_reg_0,
    D,
    \FSM_sequential_fifo_state_reg[0] ,
    \qvRAddr_reg[6]_0 ,
    \qvWAddr_reg[5]_0 ,
    fifo_rd_en,
    qEmpty_reg_1,
    qFull_reg_0,
    qFull_reg_1,
    \qvRAddr_reg[6]_1 ,
    receiving_d2,
    Q,
    \pad_cnt_reg_reg[0] ,
    fifo_rd_en_reg,
    \pad_rxc_reg_reg[0] ,
    fifo_rd_en_reg_0,
    pad_frame_d1_reg,
    clk_i,
    reset_dcm);
  output qEmpty_reg_0;
  output [2:0]D;
  output \FSM_sequential_fifo_state_reg[0] ;
  output [6:0]\qvRAddr_reg[6]_0 ;
  output [5:0]\qvWAddr_reg[5]_0 ;
  output fifo_rd_en;
  output qEmpty_reg_1;
  output qFull_reg_0;
  output qFull_reg_1;
  input \qvRAddr_reg[6]_1 ;
  input receiving_d2;
  input [2:0]Q;
  input [2:0]\pad_cnt_reg_reg[0] ;
  input [1:0]fifo_rd_en_reg;
  input \pad_rxc_reg_reg[0] ;
  input fifo_rd_en_reg_0;
  input pad_frame_d1_reg;
  input clk_i;
  input reset_dcm;

  wire [2:0]D;
  wire \FSM_sequential_fifo_state_reg[0] ;
  wire MemREn;
  wire MemWEn;
  wire [2:0]Q;
  wire clk_i;
  wire fifo_rd_en;
  wire [1:0]fifo_rd_en_reg;
  wire fifo_rd_en_reg_0;
  wire [6:0]p_0_in__0;
  wire [6:0]p_0_in__1;
  wire [2:0]\pad_cnt_reg_reg[0] ;
  wire pad_frame_d1_reg;
  wire \pad_rxc_reg_reg[0] ;
  wire qEmpty_i_1_n_0;
  wire qEmpty_i_2_n_0;
  wire qEmpty_i_3_n_0;
  wire qEmpty_reg_0;
  wire qEmpty_reg_1;
  wire qFull_i_1_n_0;
  wire qFull_i_2_n_0;
  wire qFull_i_3_n_0;
  wire qFull_reg_0;
  wire qFull_reg_1;
  wire qFull_reg_n_0;
  wire \qvCount[0]_i_1_n_0 ;
  wire \qvCount[7]_i_10_n_0 ;
  wire \qvCount[7]_i_1_n_0 ;
  wire \qvCount[7]_i_3_n_0 ;
  wire \qvCount[7]_i_4_n_0 ;
  wire \qvCount[7]_i_5_n_0 ;
  wire \qvCount[7]_i_6__0_n_0 ;
  wire \qvCount[7]_i_7_n_0 ;
  wire \qvCount[7]_i_8_n_0 ;
  wire \qvCount[7]_i_9_n_0 ;
  wire [7:0]qvCount_reg;
  wire \qvCount_reg[7]_i_2_n_10 ;
  wire \qvCount_reg[7]_i_2_n_11 ;
  wire \qvCount_reg[7]_i_2_n_12 ;
  wire \qvCount_reg[7]_i_2_n_13 ;
  wire \qvCount_reg[7]_i_2_n_14 ;
  wire \qvCount_reg[7]_i_2_n_15 ;
  wire \qvCount_reg[7]_i_2_n_2 ;
  wire \qvCount_reg[7]_i_2_n_3 ;
  wire \qvCount_reg[7]_i_2_n_4 ;
  wire \qvCount_reg[7]_i_2_n_5 ;
  wire \qvCount_reg[7]_i_2_n_6 ;
  wire \qvCount_reg[7]_i_2_n_7 ;
  wire \qvCount_reg[7]_i_2_n_9 ;
  wire \qvRAddr[6]_i_3_n_0 ;
  wire [6:0]\qvRAddr_reg[6]_0 ;
  wire \qvRAddr_reg[6]_1 ;
  wire [6:6]qvWAddr;
  wire \qvWAddr[6]_i_3_n_0 ;
  wire [5:0]\qvWAddr_reg[5]_0 ;
  wire receiving_d2;
  wire reset_dcm;
  wire [7:6]\NLW_qvCount_reg[7]_i_2_CO_UNCONNECTED ;
  wire [7:7]\NLW_qvCount_reg[7]_i_2_O_UNCONNECTED ;

  LUT4 #(
    .INIT(16'h1F00)) 
    fifo_rd_en_i_1
       (.I0(fifo_rd_en_reg[1]),
        .I1(qEmpty_reg_0),
        .I2(fifo_rd_en_reg_0),
        .I3(fifo_rd_en_reg[0]),
        .O(fifo_rd_en));
  LUT3 #(
    .INIT(8'h04)) 
    mem_reg_0_63_0_6_i_1
       (.I0(qFull_reg_n_0),
        .I1(receiving_d2),
        .I2(qvWAddr),
        .O(qFull_reg_0));
  LUT3 #(
    .INIT(8'h40)) 
    mem_reg_64_127_0_6_i_1
       (.I0(qFull_reg_n_0),
        .I1(receiving_d2),
        .I2(qvWAddr),
        .O(qFull_reg_1));
  LUT6 #(
    .INIT(64'h8B888B888B888888)) 
    \pad_cnt_reg[0]_i_1 
       (.I0(Q[0]),
        .I1(\FSM_sequential_fifo_state_reg[0] ),
        .I2(\pad_cnt_reg_reg[0] [0]),
        .I3(fifo_rd_en_reg[1]),
        .I4(\pad_cnt_reg_reg[0] [1]),
        .I5(\pad_cnt_reg_reg[0] [2]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'hB8888B88B8888888)) 
    \pad_cnt_reg[1]_i_1 
       (.I0(Q[1]),
        .I1(\FSM_sequential_fifo_state_reg[0] ),
        .I2(\pad_cnt_reg_reg[0] [0]),
        .I3(fifo_rd_en_reg[1]),
        .I4(\pad_cnt_reg_reg[0] [1]),
        .I5(\pad_cnt_reg_reg[0] [2]),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hBBB8888888888888)) 
    \pad_cnt_reg[2]_i_1 
       (.I0(Q[2]),
        .I1(\FSM_sequential_fifo_state_reg[0] ),
        .I2(\pad_cnt_reg_reg[0] [0]),
        .I3(\pad_cnt_reg_reg[0] [1]),
        .I4(\pad_cnt_reg_reg[0] [2]),
        .I5(fifo_rd_en_reg[1]),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT5 #(
    .INIT(32'hFFF00040)) 
    pad_frame_d1_i_1
       (.I0(qEmpty_reg_0),
        .I1(\pad_rxc_reg_reg[0] ),
        .I2(fifo_rd_en_reg[1]),
        .I3(fifo_rd_en_reg[0]),
        .I4(pad_frame_d1_reg),
        .O(qEmpty_reg_1));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \pad_rxc_reg[6]_i_1 
       (.I0(fifo_rd_en_reg[0]),
        .I1(fifo_rd_en_reg[1]),
        .I2(\pad_rxc_reg_reg[0] ),
        .I3(qEmpty_reg_0),
        .O(\FSM_sequential_fifo_state_reg[0] ));
  LUT6 #(
    .INIT(64'hF1F00000F1F0F1F0)) 
    qEmpty_i_1
       (.I0(qEmpty_i_2_n_0),
        .I1(qEmpty_i_3_n_0),
        .I2(qEmpty_reg_0),
        .I3(\qvRAddr_reg[6]_1 ),
        .I4(qFull_reg_n_0),
        .I5(receiving_d2),
        .O(qEmpty_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    qEmpty_i_2
       (.I0(qvCount_reg[5]),
        .I1(qvCount_reg[1]),
        .I2(qvCount_reg[0]),
        .I3(qvCount_reg[4]),
        .O(qEmpty_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    qEmpty_i_3
       (.I0(qvCount_reg[7]),
        .I1(qvCount_reg[6]),
        .I2(qvCount_reg[3]),
        .I3(qvCount_reg[2]),
        .O(qEmpty_i_3_n_0));
  FDPE #(
    .INIT(1'b1)) 
    qEmpty_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(qEmpty_i_1_n_0),
        .PRE(reset_dcm),
        .Q(qEmpty_reg_0));
  LUT6 #(
    .INIT(64'hF1F00000F1F0F1F0)) 
    qFull_i_1
       (.I0(qFull_i_2_n_0),
        .I1(qFull_i_3_n_0),
        .I2(qFull_reg_n_0),
        .I3(receiving_d2),
        .I4(qEmpty_reg_0),
        .I5(\qvRAddr_reg[6]_1 ),
        .O(qFull_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    qFull_i_2
       (.I0(qvCount_reg[6]),
        .I1(qvCount_reg[5]),
        .I2(qvCount_reg[4]),
        .O(qFull_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    qFull_i_3
       (.I0(qvCount_reg[0]),
        .I1(qvCount_reg[2]),
        .I2(qvCount_reg[3]),
        .I3(qvCount_reg[1]),
        .O(qFull_i_3_n_0));
  FDCE #(
    .INIT(1'b0)) 
    qFull_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qFull_i_1_n_0),
        .Q(qFull_reg_n_0));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \qvCount[0]_i_1 
       (.I0(qvCount_reg[0]),
        .O(\qvCount[0]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h4B44)) 
    \qvCount[7]_i_1 
       (.I0(qEmpty_reg_0),
        .I1(\qvRAddr_reg[6]_1 ),
        .I2(qFull_reg_n_0),
        .I3(receiving_d2),
        .O(\qvCount[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h65)) 
    \qvCount[7]_i_10 
       (.I0(qvCount_reg[1]),
        .I1(qFull_reg_n_0),
        .I2(receiving_d2),
        .O(\qvCount[7]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \qvCount[7]_i_3 
       (.I0(receiving_d2),
        .I1(qFull_reg_n_0),
        .O(\qvCount[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_4 
       (.I0(qvCount_reg[6]),
        .I1(qvCount_reg[7]),
        .O(\qvCount[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_5 
       (.I0(qvCount_reg[5]),
        .I1(qvCount_reg[6]),
        .O(\qvCount[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_6__0 
       (.I0(qvCount_reg[4]),
        .I1(qvCount_reg[5]),
        .O(\qvCount[7]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_7 
       (.I0(qvCount_reg[3]),
        .I1(qvCount_reg[4]),
        .O(\qvCount[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_8 
       (.I0(qvCount_reg[2]),
        .I1(qvCount_reg[3]),
        .O(\qvCount[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_9 
       (.I0(qvCount_reg[1]),
        .I1(qvCount_reg[2]),
        .O(\qvCount[7]_i_9_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[0] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount[0]_i_1_n_0 ),
        .Q(qvCount_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[1] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_15 ),
        .Q(qvCount_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[2] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_14 ),
        .Q(qvCount_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[3] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_13 ),
        .Q(qvCount_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[4] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_12 ),
        .Q(qvCount_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[5] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_11 ),
        .Q(qvCount_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[6] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_10 ),
        .Q(qvCount_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[7] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2_n_9 ),
        .Q(qvCount_reg[7]));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \qvCount_reg[7]_i_2 
       (.CI(qvCount_reg[0]),
        .CI_TOP(1'b0),
        .CO({\NLW_qvCount_reg[7]_i_2_CO_UNCONNECTED [7:6],\qvCount_reg[7]_i_2_n_2 ,\qvCount_reg[7]_i_2_n_3 ,\qvCount_reg[7]_i_2_n_4 ,\qvCount_reg[7]_i_2_n_5 ,\qvCount_reg[7]_i_2_n_6 ,\qvCount_reg[7]_i_2_n_7 }),
        .DI({1'b0,1'b0,qvCount_reg[5:1],\qvCount[7]_i_3_n_0 }),
        .O({\NLW_qvCount_reg[7]_i_2_O_UNCONNECTED [7],\qvCount_reg[7]_i_2_n_9 ,\qvCount_reg[7]_i_2_n_10 ,\qvCount_reg[7]_i_2_n_11 ,\qvCount_reg[7]_i_2_n_12 ,\qvCount_reg[7]_i_2_n_13 ,\qvCount_reg[7]_i_2_n_14 ,\qvCount_reg[7]_i_2_n_15 }),
        .S({1'b0,\qvCount[7]_i_4_n_0 ,\qvCount[7]_i_5_n_0 ,\qvCount[7]_i_6__0_n_0 ,\qvCount[7]_i_7_n_0 ,\qvCount[7]_i_8_n_0 ,\qvCount[7]_i_9_n_0 ,\qvCount[7]_i_10_n_0 }));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \qvRAddr[0]_i_1 
       (.I0(\qvRAddr_reg[6]_0 [0]),
        .O(p_0_in__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRAddr[1]_i_1 
       (.I0(\qvRAddr_reg[6]_0 [0]),
        .I1(\qvRAddr_reg[6]_0 [1]),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \qvRAddr[2]_i_1 
       (.I0(\qvRAddr_reg[6]_0 [2]),
        .I1(\qvRAddr_reg[6]_0 [0]),
        .I2(\qvRAddr_reg[6]_0 [1]),
        .O(p_0_in__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \qvRAddr[3]_i_1 
       (.I0(\qvRAddr_reg[6]_0 [3]),
        .I1(\qvRAddr_reg[6]_0 [1]),
        .I2(\qvRAddr_reg[6]_0 [0]),
        .I3(\qvRAddr_reg[6]_0 [2]),
        .O(p_0_in__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \qvRAddr[4]_i_1 
       (.I0(\qvRAddr_reg[6]_0 [4]),
        .I1(\qvRAddr_reg[6]_0 [2]),
        .I2(\qvRAddr_reg[6]_0 [0]),
        .I3(\qvRAddr_reg[6]_0 [1]),
        .I4(\qvRAddr_reg[6]_0 [3]),
        .O(p_0_in__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \qvRAddr[5]_i_1 
       (.I0(\qvRAddr_reg[6]_0 [3]),
        .I1(\qvRAddr_reg[6]_0 [1]),
        .I2(\qvRAddr_reg[6]_0 [0]),
        .I3(\qvRAddr_reg[6]_0 [2]),
        .I4(\qvRAddr_reg[6]_0 [4]),
        .I5(\qvRAddr_reg[6]_0 [5]),
        .O(p_0_in__0[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \qvRAddr[6]_i_1 
       (.I0(\qvRAddr_reg[6]_1 ),
        .I1(qEmpty_reg_0),
        .O(MemREn));
  LUT3 #(
    .INIT(8'h9A)) 
    \qvRAddr[6]_i_2 
       (.I0(\qvRAddr_reg[6]_0 [6]),
        .I1(\qvRAddr[6]_i_3_n_0 ),
        .I2(\qvRAddr_reg[6]_0 [5]),
        .O(p_0_in__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \qvRAddr[6]_i_3 
       (.I0(\qvRAddr_reg[6]_0 [3]),
        .I1(\qvRAddr_reg[6]_0 [1]),
        .I2(\qvRAddr_reg[6]_0 [0]),
        .I3(\qvRAddr_reg[6]_0 [2]),
        .I4(\qvRAddr_reg[6]_0 [4]),
        .O(\qvRAddr[6]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[0] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[0]),
        .Q(\qvRAddr_reg[6]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[1] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[1]),
        .Q(\qvRAddr_reg[6]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[2] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[2]),
        .Q(\qvRAddr_reg[6]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[3] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[3]),
        .Q(\qvRAddr_reg[6]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[4] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[4]),
        .Q(\qvRAddr_reg[6]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[5] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[5]),
        .Q(\qvRAddr_reg[6]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[6] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__0[6]),
        .Q(\qvRAddr_reg[6]_0 [6]));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \qvWAddr[0]_i_1 
       (.I0(\qvWAddr_reg[5]_0 [0]),
        .O(p_0_in__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvWAddr[1]_i_1 
       (.I0(\qvWAddr_reg[5]_0 [0]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .O(p_0_in__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \qvWAddr[2]_i_1 
       (.I0(\qvWAddr_reg[5]_0 [2]),
        .I1(\qvWAddr_reg[5]_0 [0]),
        .I2(\qvWAddr_reg[5]_0 [1]),
        .O(p_0_in__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \qvWAddr[3]_i_1 
       (.I0(\qvWAddr_reg[5]_0 [3]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [2]),
        .O(p_0_in__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \qvWAddr[4]_i_1__0 
       (.I0(\qvWAddr_reg[5]_0 [4]),
        .I1(\qvWAddr_reg[5]_0 [2]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [1]),
        .I4(\qvWAddr_reg[5]_0 [3]),
        .O(p_0_in__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \qvWAddr[5]_i_1 
       (.I0(\qvWAddr_reg[5]_0 [3]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [2]),
        .I4(\qvWAddr_reg[5]_0 [4]),
        .I5(\qvWAddr_reg[5]_0 [5]),
        .O(p_0_in__1[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \qvWAddr[6]_i_1 
       (.I0(receiving_d2),
        .I1(qFull_reg_n_0),
        .O(MemWEn));
  LUT3 #(
    .INIT(8'h9A)) 
    \qvWAddr[6]_i_2 
       (.I0(qvWAddr),
        .I1(\qvWAddr[6]_i_3_n_0 ),
        .I2(\qvWAddr_reg[5]_0 [5]),
        .O(p_0_in__1[6]));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \qvWAddr[6]_i_3 
       (.I0(\qvWAddr_reg[5]_0 [3]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [2]),
        .I4(\qvWAddr_reg[5]_0 [4]),
        .O(\qvWAddr[6]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[0] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[0]),
        .Q(\qvWAddr_reg[5]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[1] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[1]),
        .Q(\qvWAddr_reg[5]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[2] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[2]),
        .Q(\qvWAddr_reg[5]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[3] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[3]),
        .Q(\qvWAddr_reg[5]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[4] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[4]),
        .Q(\qvWAddr_reg[5]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[5] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[5]),
        .Q(\qvWAddr_reg[5]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[6] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__1[6]),
        .Q(qvWAddr));
endmodule

(* ORIG_REF_NAME = "FifoControl" *) 
module switch_elements_FifoControl_2
   (qEmpty_reg_0,
    Q,
    \qvWAddr_reg[5]_0 ,
    qFull_reg_0,
    qFull_reg_1,
    \qvRAddr_reg[6]_0 ,
    receiving_d2,
    clk_i,
    reset_dcm);
  output qEmpty_reg_0;
  output [6:0]Q;
  output [5:0]\qvWAddr_reg[5]_0 ;
  output qFull_reg_0;
  output qFull_reg_1;
  input \qvRAddr_reg[6]_0 ;
  input receiving_d2;
  input clk_i;
  input reset_dcm;

  wire MemREn;
  wire MemWEn;
  wire [6:0]Q;
  wire clk_i;
  wire [6:0]p_0_in__3;
  wire [6:0]p_0_in__4;
  wire qEmpty_i_1_n_0;
  wire qEmpty_i_2__0_n_0;
  wire qEmpty_i_3__0_n_0;
  wire qEmpty_reg_0;
  wire qFull_i_1_n_0;
  wire qFull_i_2__0_n_0;
  wire qFull_i_3__0_n_0;
  wire qFull_reg_0;
  wire qFull_reg_1;
  wire qFull_reg_n_0;
  wire \qvCount[0]_i_1__0_n_0 ;
  wire \qvCount[7]_i_10__0_n_0 ;
  wire \qvCount[7]_i_1__0_n_0 ;
  wire \qvCount[7]_i_3__0_n_0 ;
  wire \qvCount[7]_i_4__0_n_0 ;
  wire \qvCount[7]_i_5__0_n_0 ;
  wire \qvCount[7]_i_6_n_0 ;
  wire \qvCount[7]_i_7__0_n_0 ;
  wire \qvCount[7]_i_8__0_n_0 ;
  wire \qvCount[7]_i_9__0_n_0 ;
  wire [7:0]qvCount_reg;
  wire \qvCount_reg[7]_i_2__0_n_10 ;
  wire \qvCount_reg[7]_i_2__0_n_11 ;
  wire \qvCount_reg[7]_i_2__0_n_12 ;
  wire \qvCount_reg[7]_i_2__0_n_13 ;
  wire \qvCount_reg[7]_i_2__0_n_14 ;
  wire \qvCount_reg[7]_i_2__0_n_15 ;
  wire \qvCount_reg[7]_i_2__0_n_2 ;
  wire \qvCount_reg[7]_i_2__0_n_3 ;
  wire \qvCount_reg[7]_i_2__0_n_4 ;
  wire \qvCount_reg[7]_i_2__0_n_5 ;
  wire \qvCount_reg[7]_i_2__0_n_6 ;
  wire \qvCount_reg[7]_i_2__0_n_7 ;
  wire \qvCount_reg[7]_i_2__0_n_9 ;
  wire \qvRAddr[6]_i_3__0_n_0 ;
  wire \qvRAddr_reg[6]_0 ;
  wire \qvWAddr[6]_i_3__0_n_0 ;
  wire [5:0]\qvWAddr_reg[5]_0 ;
  wire \qvWAddr_reg_n_0_[6] ;
  wire receiving_d2;
  wire reset_dcm;
  wire [7:6]\NLW_qvCount_reg[7]_i_2__0_CO_UNCONNECTED ;
  wire [7:7]\NLW_qvCount_reg[7]_i_2__0_O_UNCONNECTED ;

  LUT3 #(
    .INIT(8'h04)) 
    mem_reg_0_63_0_6_i_8
       (.I0(qFull_reg_n_0),
        .I1(receiving_d2),
        .I2(\qvWAddr_reg_n_0_[6] ),
        .O(qFull_reg_0));
  LUT3 #(
    .INIT(8'h40)) 
    mem_reg_64_127_0_6_i_1__0
       (.I0(qFull_reg_n_0),
        .I1(receiving_d2),
        .I2(\qvWAddr_reg_n_0_[6] ),
        .O(qFull_reg_1));
  LUT6 #(
    .INIT(64'hF1F00000F1F0F1F0)) 
    qEmpty_i_1
       (.I0(qEmpty_i_2__0_n_0),
        .I1(qEmpty_i_3__0_n_0),
        .I2(qEmpty_reg_0),
        .I3(\qvRAddr_reg[6]_0 ),
        .I4(qFull_reg_n_0),
        .I5(receiving_d2),
        .O(qEmpty_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    qEmpty_i_2__0
       (.I0(qvCount_reg[0]),
        .I1(qvCount_reg[1]),
        .I2(qvCount_reg[5]),
        .I3(qvCount_reg[4]),
        .O(qEmpty_i_2__0_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    qEmpty_i_3__0
       (.I0(qvCount_reg[7]),
        .I1(qvCount_reg[6]),
        .I2(qvCount_reg[3]),
        .I3(qvCount_reg[2]),
        .O(qEmpty_i_3__0_n_0));
  FDPE #(
    .INIT(1'b1)) 
    qEmpty_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(qEmpty_i_1_n_0),
        .PRE(reset_dcm),
        .Q(qEmpty_reg_0));
  LUT6 #(
    .INIT(64'hF1F00000F1F0F1F0)) 
    qFull_i_1
       (.I0(qFull_i_2__0_n_0),
        .I1(qFull_i_3__0_n_0),
        .I2(qFull_reg_n_0),
        .I3(receiving_d2),
        .I4(qEmpty_reg_0),
        .I5(\qvRAddr_reg[6]_0 ),
        .O(qFull_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    qFull_i_2__0
       (.I0(qvCount_reg[6]),
        .I1(qvCount_reg[1]),
        .I2(qvCount_reg[5]),
        .O(qFull_i_2__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    qFull_i_3__0
       (.I0(qvCount_reg[4]),
        .I1(qvCount_reg[3]),
        .I2(qvCount_reg[0]),
        .I3(qvCount_reg[2]),
        .O(qFull_i_3__0_n_0));
  FDCE #(
    .INIT(1'b0)) 
    qFull_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qFull_i_1_n_0),
        .Q(qFull_reg_n_0));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \qvCount[0]_i_1__0 
       (.I0(qvCount_reg[0]),
        .O(\qvCount[0]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'h65)) 
    \qvCount[7]_i_10__0 
       (.I0(qvCount_reg[1]),
        .I1(qFull_reg_n_0),
        .I2(receiving_d2),
        .O(\qvCount[7]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h4B44)) 
    \qvCount[7]_i_1__0 
       (.I0(qEmpty_reg_0),
        .I1(\qvRAddr_reg[6]_0 ),
        .I2(qFull_reg_n_0),
        .I3(receiving_d2),
        .O(\qvCount[7]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \qvCount[7]_i_3__0 
       (.I0(receiving_d2),
        .I1(qFull_reg_n_0),
        .O(\qvCount[7]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_4__0 
       (.I0(qvCount_reg[6]),
        .I1(qvCount_reg[7]),
        .O(\qvCount[7]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_5__0 
       (.I0(qvCount_reg[5]),
        .I1(qvCount_reg[6]),
        .O(\qvCount[7]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_6 
       (.I0(qvCount_reg[4]),
        .I1(qvCount_reg[5]),
        .O(\qvCount[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_7__0 
       (.I0(qvCount_reg[3]),
        .I1(qvCount_reg[4]),
        .O(\qvCount[7]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_8__0 
       (.I0(qvCount_reg[2]),
        .I1(qvCount_reg[3]),
        .O(\qvCount[7]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \qvCount[7]_i_9__0 
       (.I0(qvCount_reg[1]),
        .I1(qvCount_reg[2]),
        .O(\qvCount[7]_i_9__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[0] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount[0]_i_1__0_n_0 ),
        .Q(qvCount_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[1] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_15 ),
        .Q(qvCount_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[2] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_14 ),
        .Q(qvCount_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[3] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_13 ),
        .Q(qvCount_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[4] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_12 ),
        .Q(qvCount_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[5] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_11 ),
        .Q(qvCount_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[6] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_10 ),
        .Q(qvCount_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \qvCount_reg[7] 
       (.C(clk_i),
        .CE(\qvCount[7]_i_1__0_n_0 ),
        .CLR(reset_dcm),
        .D(\qvCount_reg[7]_i_2__0_n_9 ),
        .Q(qvCount_reg[7]));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \qvCount_reg[7]_i_2__0 
       (.CI(qvCount_reg[0]),
        .CI_TOP(1'b0),
        .CO({\NLW_qvCount_reg[7]_i_2__0_CO_UNCONNECTED [7:6],\qvCount_reg[7]_i_2__0_n_2 ,\qvCount_reg[7]_i_2__0_n_3 ,\qvCount_reg[7]_i_2__0_n_4 ,\qvCount_reg[7]_i_2__0_n_5 ,\qvCount_reg[7]_i_2__0_n_6 ,\qvCount_reg[7]_i_2__0_n_7 }),
        .DI({1'b0,1'b0,qvCount_reg[5:1],\qvCount[7]_i_3__0_n_0 }),
        .O({\NLW_qvCount_reg[7]_i_2__0_O_UNCONNECTED [7],\qvCount_reg[7]_i_2__0_n_9 ,\qvCount_reg[7]_i_2__0_n_10 ,\qvCount_reg[7]_i_2__0_n_11 ,\qvCount_reg[7]_i_2__0_n_12 ,\qvCount_reg[7]_i_2__0_n_13 ,\qvCount_reg[7]_i_2__0_n_14 ,\qvCount_reg[7]_i_2__0_n_15 }),
        .S({1'b0,\qvCount[7]_i_4__0_n_0 ,\qvCount[7]_i_5__0_n_0 ,\qvCount[7]_i_6_n_0 ,\qvCount[7]_i_7__0_n_0 ,\qvCount[7]_i_8__0_n_0 ,\qvCount[7]_i_9__0_n_0 ,\qvCount[7]_i_10__0_n_0 }));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \qvRAddr[0]_i_1__0 
       (.I0(Q[0]),
        .O(p_0_in__3[0]));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRAddr[1]_i_1__0 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(p_0_in__3[1]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \qvRAddr[2]_i_1__0 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(p_0_in__3[2]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \qvRAddr[3]_i_1__0 
       (.I0(Q[3]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[2]),
        .O(p_0_in__3[3]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \qvRAddr[4]_i_1__0 
       (.I0(Q[4]),
        .I1(Q[2]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(Q[3]),
        .O(p_0_in__3[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \qvRAddr[5]_i_1__0 
       (.I0(Q[3]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(Q[4]),
        .I5(Q[5]),
        .O(p_0_in__3[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \qvRAddr[6]_i_1__0 
       (.I0(\qvRAddr_reg[6]_0 ),
        .I1(qEmpty_reg_0),
        .O(MemREn));
  LUT3 #(
    .INIT(8'h9A)) 
    \qvRAddr[6]_i_2__0 
       (.I0(Q[6]),
        .I1(\qvRAddr[6]_i_3__0_n_0 ),
        .I2(Q[5]),
        .O(p_0_in__3[6]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \qvRAddr[6]_i_3__0 
       (.I0(Q[3]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(Q[4]),
        .O(\qvRAddr[6]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[0] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[0]),
        .Q(Q[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[1] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[1]),
        .Q(Q[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[2] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[2]),
        .Q(Q[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[3] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[3]),
        .Q(Q[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[4] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[4]),
        .Q(Q[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[5] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[5]),
        .Q(Q[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[6] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(reset_dcm),
        .D(p_0_in__3[6]),
        .Q(Q[6]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \qvWAddr[0]_i_1__0 
       (.I0(\qvWAddr_reg[5]_0 [0]),
        .O(p_0_in__4[0]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvWAddr[1]_i_1__0 
       (.I0(\qvWAddr_reg[5]_0 [0]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .O(p_0_in__4[1]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \qvWAddr[2]_i_1__0 
       (.I0(\qvWAddr_reg[5]_0 [2]),
        .I1(\qvWAddr_reg[5]_0 [0]),
        .I2(\qvWAddr_reg[5]_0 [1]),
        .O(p_0_in__4[2]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \qvWAddr[3]_i_1__0 
       (.I0(\qvWAddr_reg[5]_0 [3]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [2]),
        .O(p_0_in__4[3]));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \qvWAddr[4]_i_1__1 
       (.I0(\qvWAddr_reg[5]_0 [4]),
        .I1(\qvWAddr_reg[5]_0 [2]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [1]),
        .I4(\qvWAddr_reg[5]_0 [3]),
        .O(p_0_in__4[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \qvWAddr[5]_i_1__0 
       (.I0(\qvWAddr_reg[5]_0 [3]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [2]),
        .I4(\qvWAddr_reg[5]_0 [4]),
        .I5(\qvWAddr_reg[5]_0 [5]),
        .O(p_0_in__4[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \qvWAddr[6]_i_1__0 
       (.I0(receiving_d2),
        .I1(qFull_reg_n_0),
        .O(MemWEn));
  LUT3 #(
    .INIT(8'h9A)) 
    \qvWAddr[6]_i_2__0 
       (.I0(\qvWAddr_reg_n_0_[6] ),
        .I1(\qvWAddr[6]_i_3__0_n_0 ),
        .I2(\qvWAddr_reg[5]_0 [5]),
        .O(p_0_in__4[6]));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \qvWAddr[6]_i_3__0 
       (.I0(\qvWAddr_reg[5]_0 [3]),
        .I1(\qvWAddr_reg[5]_0 [1]),
        .I2(\qvWAddr_reg[5]_0 [0]),
        .I3(\qvWAddr_reg[5]_0 [2]),
        .I4(\qvWAddr_reg[5]_0 [4]),
        .O(\qvWAddr[6]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[0] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[0]),
        .Q(\qvWAddr_reg[5]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[1] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[1]),
        .Q(\qvWAddr_reg[5]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[2] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[2]),
        .Q(\qvWAddr_reg[5]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[3] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[3]),
        .Q(\qvWAddr_reg[5]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[4] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[4]),
        .Q(\qvWAddr_reg[5]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[5] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[5]),
        .Q(\qvWAddr_reg[5]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[6] 
       (.C(clk_i),
        .CE(MemWEn),
        .CLR(reset_dcm),
        .D(p_0_in__4[6]),
        .Q(\qvWAddr_reg_n_0_[6] ));
endmodule

(* ORIG_REF_NAME = "FifoControl_ASYN" *) 
module switch_elements_FifoControl_ASYN
   (rst_i_0,
    ADDRH,
    E,
    D,
    this_cycle,
    \qvDataOut_reg[25]_0 ,
    \qvDataOut_reg[66]_0 ,
    \qvDataOut_reg[71]_0 ,
    \qvDataOut_reg[69]_0 ,
    \qvDataOut_reg[62]_0 ,
    get_sfd0,
    \qvDataOut_reg[45]_0 ,
    clk_i,
    Q,
    \qvDataOut_reg[71]_1 ,
    rst_i,
    recv_rst);
  output rst_i_0;
  output [4:0]ADDRH;
  output [0:0]E;
  output [4:0]D;
  output this_cycle;
  output [5:0]\qvDataOut_reg[25]_0 ;
  output [0:0]\qvDataOut_reg[66]_0 ;
  output [71:0]\qvDataOut_reg[71]_0 ;
  output [2:0]\qvDataOut_reg[69]_0 ;
  output [7:0]\qvDataOut_reg[62]_0 ;
  output get_sfd0;
  output \qvDataOut_reg[45]_0 ;
  input clk_i;
  input [0:0]Q;
  input [71:0]\qvDataOut_reg[71]_1 ;
  input rst_i;
  input recv_rst;

  wire [4:0]ADDRH;
  wire [4:0]D;
  wire [0:0]E;
  wire MemREn;
  wire [0:0]Q;
  wire \_inferred__1/i__carry_n_3 ;
  wire \_inferred__1/i__carry_n_4 ;
  wire \_inferred__1/i__carry_n_5 ;
  wire \_inferred__1/i__carry_n_6 ;
  wire \_inferred__1/i__carry_n_7 ;
  wire clk_i;
  wire \get_e_chk[0]_i_2_n_0 ;
  wire \get_e_chk[1]_i_2_n_0 ;
  wire \get_e_chk[2]_i_2_n_0 ;
  wire \get_e_chk[3]_i_2_n_0 ;
  wire \get_e_chk[4]_i_2_n_0 ;
  wire \get_e_chk[5]_i_2_n_0 ;
  wire \get_e_chk[6]_i_2_n_0 ;
  wire \get_e_chk[7]_i_2_n_0 ;
  wire get_sfd0;
  wire get_sfd_i_2_n_0;
  wire get_sfd_i_3_n_0;
  wire get_sfd_i_4_n_0;
  wire get_sfd_i_5_n_0;
  wire i__carry_i_10__3_n_0;
  wire i__carry_i_11_n_0;
  wire i__carry_i_1__3_n_0;
  wire i__carry_i_2__3_n_0;
  wire i__carry_i_3__3_n_0;
  wire i__carry_i_4__3_n_0;
  wire i__carry_i_5__3_n_0;
  wire i__carry_i_6__2_n_0;
  wire i__carry_i_7__2_n_0;
  wire i__carry_i_8__1_n_0;
  wire i__carry_i_9__2_n_0;
  wire [5:0]p_0_in__2;
  wire [5:0]p_0_in__5;
  wire qREmpty_int_i_1_n_0;
  wire qREmpty_int_i_2_n_0;
  wire qREmpty_int_i_3_n_0;
  wire qREmpty_int_i_4_n_0;
  wire qREmpty_int_i_5_n_0;
  wire qREmpty_int_reg_n_0;
  wire [5:0]\qvDataOut_reg[25]_0 ;
  wire \qvDataOut_reg[45]_0 ;
  wire [7:0]\qvDataOut_reg[62]_0 ;
  wire [0:0]\qvDataOut_reg[66]_0 ;
  wire [2:0]\qvDataOut_reg[69]_0 ;
  wire [71:0]\qvDataOut_reg[71]_0 ;
  wire [71:0]\qvDataOut_reg[71]_1 ;
  wire [5:0]qvNextRAddr_reg;
  wire [5:0]qvNextWAddr_reg;
  wire [5:1]qvPreWGrayAddr;
  wire [5:0]qvPreWGrayAddr_RSync1;
  wire [5:0]qvPreWGrayAddr_RSync2;
  wire [4:0]qvRAddr;
  wire [5:0]qvRAddr_WSync2;
  wire qvRAddr_WSync20__0;
  wire \qvRAddr_WSync20_inferred__0/i__n_0 ;
  wire qvRAddr_WSync20_n_0;
  wire \qvRAddr_WSync2[2]_i_1_n_0 ;
  wire \qvRAddr_WSync2[3]_i_1_n_0 ;
  wire [5:0]qvRGrayAddr;
  wire [4:0]qvRGrayAddr0;
  wire [5:0]qvRGrayAddr_WSync1;
  wire [5:0]qvRGrayAddr_WSync2;
  wire [5:5]qvWCount;
  wire \qvWCount_reg_n_0_[5] ;
  wire [4:1]qvWGrayAddr;
  wire [4:0]qvWGrayAddr0;
  wire [5:0]qvWGrayAddr_RSync1;
  wire [5:0]qvWGrayAddr_RSync2;
  wire recv_rst;
  wire rst_i;
  wire rst_i_0;
  wire \rxc_end_data[2]_i_2_n_0 ;
  wire \rxc_end_data[4]_i_2_n_0 ;
  wire \rxc_end_data[4]_i_3_n_0 ;
  wire \rxc_end_data[4]_i_4_n_0 ;
  wire \rxc_end_data[7]_i_10_n_0 ;
  wire \rxc_end_data[7]_i_3_n_0 ;
  wire \rxc_end_data[7]_i_4_n_0 ;
  wire \rxc_end_data[7]_i_5_n_0 ;
  wire \rxc_end_data[7]_i_6_n_0 ;
  wire \rxc_end_data[7]_i_7_n_0 ;
  wire \rxc_end_data[7]_i_8_n_0 ;
  wire \rxc_end_data[7]_i_9_n_0 ;
  wire tagged_frame_i_2_n_0;
  wire tagged_frame_i_3_n_0;
  wire tagged_frame_i_4_n_0;
  wire tagged_frame_i_5_n_0;
  wire tagged_frame_i_6_n_0;
  wire tagged_frame_i_7_n_0;
  wire tagged_frame_i_8_n_0;
  wire tagged_frame_i_9_n_0;
  wire \terminator_location[0]_i_2_n_0 ;
  wire \terminator_location[0]_i_3_n_0 ;
  wire \terminator_location[0]_i_4_n_0 ;
  wire \terminator_location[1]_i_2_n_0 ;
  wire \terminator_location[1]_i_3_n_0 ;
  wire this_cycle;
  wire [5:5]vWAddr;
  wire [7:5]\NLW__inferred__1/i__carry_CO_UNCONNECTED ;
  wire [7:0]\NLW__inferred__1/i__carry_O_UNCONNECTED ;

  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_fifo_state[1]_i_2 
       (.I0(rst_i),
        .I1(recv_rst),
        .O(rst_i_0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \_inferred__1/i__carry 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\NLW__inferred__1/i__carry_CO_UNCONNECTED [7:5],\_inferred__1/i__carry_n_3 ,\_inferred__1/i__carry_n_4 ,\_inferred__1/i__carry_n_5 ,\_inferred__1/i__carry_n_6 ,\_inferred__1/i__carry_n_7 }),
        .DI({1'b0,1'b0,1'b0,i__carry_i_1__3_n_0,i__carry_i_2__3_n_0,i__carry_i_3__3_n_0,i__carry_i_4__3_n_0,i__carry_i_5__3_n_0}),
        .O({\NLW__inferred__1/i__carry_O_UNCONNECTED [7:6],qvWCount,\NLW__inferred__1/i__carry_O_UNCONNECTED [4:0]}),
        .S({1'b0,1'b0,i__carry_i_6__2_n_0,i__carry_i_7__2_n_0,i__carry_i_8__1_n_0,i__carry_i_9__2_n_0,i__carry_i_10__3_n_0,i__carry_i_11_n_0}));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \get_e_chk[0]_i_1 
       (.I0(\qvDataOut_reg[71]_0 [0]),
        .I1(\qvDataOut_reg[71]_0 [64]),
        .I2(\qvDataOut_reg[71]_0 [3]),
        .I3(\qvDataOut_reg[71]_0 [6]),
        .I4(\qvDataOut_reg[71]_0 [2]),
        .I5(\get_e_chk[0]_i_2_n_0 ),
        .O(\qvDataOut_reg[62]_0 [0]));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \get_e_chk[0]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [5]),
        .I1(\qvDataOut_reg[71]_0 [4]),
        .I2(\qvDataOut_reg[71]_0 [7]),
        .I3(\qvDataOut_reg[71]_0 [1]),
        .O(\get_e_chk[0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT5 #(
    .INIT(32'h20000000)) 
    \get_e_chk[1]_i_1 
       (.I0(\get_e_chk[1]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [8]),
        .I2(\qvDataOut_reg[71]_0 [15]),
        .I3(\qvDataOut_reg[71]_0 [65]),
        .I4(\qvDataOut_reg[71]_0 [9]),
        .O(\qvDataOut_reg[62]_0 [1]));
  LUT5 #(
    .INIT(32'h80000000)) 
    \get_e_chk[1]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [11]),
        .I1(\qvDataOut_reg[71]_0 [10]),
        .I2(\qvDataOut_reg[71]_0 [13]),
        .I3(\qvDataOut_reg[71]_0 [14]),
        .I4(\qvDataOut_reg[71]_0 [12]),
        .O(\get_e_chk[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \get_e_chk[2]_i_1 
       (.I0(\qvDataOut_reg[71]_0 [66]),
        .I1(\get_e_chk[2]_i_2_n_0 ),
        .I2(\qvDataOut_reg[71]_0 [19]),
        .I3(\qvDataOut_reg[71]_0 [18]),
        .I4(\qvDataOut_reg[71]_0 [17]),
        .I5(\qvDataOut_reg[71]_0 [23]),
        .O(\qvDataOut_reg[62]_0 [2]));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT4 #(
    .INIT(16'hFF7F)) 
    \get_e_chk[2]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [21]),
        .I1(\qvDataOut_reg[71]_0 [20]),
        .I2(\qvDataOut_reg[71]_0 [22]),
        .I3(\qvDataOut_reg[71]_0 [16]),
        .O(\get_e_chk[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT5 #(
    .INIT(32'h20000000)) 
    \get_e_chk[3]_i_1 
       (.I0(\get_e_chk[3]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [24]),
        .I2(\qvDataOut_reg[71]_0 [25]),
        .I3(\qvDataOut_reg[71]_0 [26]),
        .I4(\qvDataOut_reg[71]_0 [27]),
        .O(\qvDataOut_reg[62]_0 [3]));
  LUT5 #(
    .INIT(32'h80000000)) 
    \get_e_chk[3]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [29]),
        .I1(\qvDataOut_reg[71]_0 [28]),
        .I2(\qvDataOut_reg[71]_0 [67]),
        .I3(\qvDataOut_reg[71]_0 [30]),
        .I4(\qvDataOut_reg[71]_0 [31]),
        .O(\get_e_chk[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \get_e_chk[4]_i_1 
       (.I0(\get_e_chk[4]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [39]),
        .I2(\qvDataOut_reg[71]_0 [32]),
        .I3(\qvDataOut_reg[71]_0 [33]),
        .I4(\qvDataOut_reg[71]_0 [68]),
        .I5(\qvDataOut_reg[71]_0 [38]),
        .O(\qvDataOut_reg[62]_0 [4]));
  LUT4 #(
    .INIT(16'h8000)) 
    \get_e_chk[4]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [37]),
        .I1(\qvDataOut_reg[71]_0 [36]),
        .I2(\qvDataOut_reg[71]_0 [35]),
        .I3(\qvDataOut_reg[71]_0 [34]),
        .O(\get_e_chk[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \get_e_chk[5]_i_1 
       (.I0(\get_e_chk[5]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [69]),
        .I2(\qvDataOut_reg[71]_0 [41]),
        .I3(\qvDataOut_reg[71]_0 [40]),
        .O(\qvDataOut_reg[62]_0 [5]));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \get_e_chk[5]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [45]),
        .I1(\qvDataOut_reg[71]_0 [43]),
        .I2(\qvDataOut_reg[71]_0 [44]),
        .I3(\qvDataOut_reg[71]_0 [46]),
        .I4(\qvDataOut_reg[71]_0 [42]),
        .I5(\qvDataOut_reg[71]_0 [47]),
        .O(\get_e_chk[5]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \get_e_chk[6]_i_1 
       (.I0(\get_e_chk[6]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [70]),
        .I2(\qvDataOut_reg[71]_0 [49]),
        .I3(\qvDataOut_reg[71]_0 [48]),
        .O(\qvDataOut_reg[62]_0 [6]));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \get_e_chk[6]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [53]),
        .I1(\qvDataOut_reg[71]_0 [51]),
        .I2(\qvDataOut_reg[71]_0 [52]),
        .I3(\qvDataOut_reg[71]_0 [54]),
        .I4(\qvDataOut_reg[71]_0 [50]),
        .I5(\qvDataOut_reg[71]_0 [55]),
        .O(\get_e_chk[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \get_e_chk[7]_i_1 
       (.I0(\qvDataOut_reg[71]_0 [62]),
        .I1(\qvDataOut_reg[71]_0 [56]),
        .I2(\qvDataOut_reg[71]_0 [57]),
        .I3(\qvDataOut_reg[71]_0 [63]),
        .I4(\qvDataOut_reg[71]_0 [71]),
        .I5(\get_e_chk[7]_i_2_n_0 ),
        .O(\qvDataOut_reg[62]_0 [7]));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \get_e_chk[7]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [59]),
        .I1(\qvDataOut_reg[71]_0 [58]),
        .I2(\qvDataOut_reg[71]_0 [61]),
        .I3(\qvDataOut_reg[71]_0 [60]),
        .O(\get_e_chk[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    get_sfd_i_1
       (.I0(get_sfd_i_2_n_0),
        .I1(\qvDataOut_reg[71]_0 [61]),
        .I2(\qvDataOut_reg[71]_0 [0]),
        .I3(\qvDataOut_reg[71]_0 [6]),
        .I4(\qvDataOut_reg[71]_0 [70]),
        .I5(get_sfd_i_3_n_0),
        .O(get_sfd0));
  LUT4 #(
    .INIT(16'hFFFD)) 
    get_sfd_i_2
       (.I0(\qvDataOut_reg[71]_0 [60]),
        .I1(\qvDataOut_reg[71]_0 [59]),
        .I2(\qvDataOut_reg[71]_0 [65]),
        .I3(\qvDataOut_reg[71]_0 [66]),
        .O(get_sfd_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    get_sfd_i_3
       (.I0(get_sfd_i_4_n_0),
        .I1(\qvDataOut_reg[71]_0 [64]),
        .I2(\qvDataOut_reg[71]_0 [69]),
        .I3(\qvDataOut_reg[71]_0 [3]),
        .I4(\qvDataOut_reg[71]_0 [67]),
        .I5(get_sfd_i_5_n_0),
        .O(get_sfd_i_3_n_0));
  LUT4 #(
    .INIT(16'hFFFD)) 
    get_sfd_i_4
       (.I0(\qvDataOut_reg[71]_0 [58]),
        .I1(\qvDataOut_reg[71]_0 [68]),
        .I2(\qvDataOut_reg[71]_0 [71]),
        .I3(\qvDataOut_reg[71]_0 [2]),
        .O(get_sfd_i_4_n_0));
  LUT5 #(
    .INIT(32'hFFFFBFFF)) 
    get_sfd_i_5
       (.I0(\qvDataOut_reg[71]_0 [57]),
        .I1(\qvDataOut_reg[71]_0 [62]),
        .I2(\qvDataOut_reg[71]_0 [56]),
        .I3(\qvDataOut_reg[71]_0 [63]),
        .I4(\get_e_chk[0]_i_2_n_0 ),
        .O(get_sfd_i_5_n_0));
  LUT5 #(
    .INIT(32'h9A999599)) 
    i__carry_i_10__3
       (.I0(qvRAddr_WSync2[1]),
        .I1(ADDRH[1]),
        .I2(\qvWCount_reg_n_0_[5] ),
        .I3(Q),
        .I4(qvNextWAddr_reg[1]),
        .O(i__carry_i_10__3_n_0));
  LUT5 #(
    .INIT(32'h9A999599)) 
    i__carry_i_11
       (.I0(qvRAddr_WSync2[0]),
        .I1(ADDRH[0]),
        .I2(\qvWCount_reg_n_0_[5] ),
        .I3(Q),
        .I4(qvNextWAddr_reg[0]),
        .O(i__carry_i_11_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_1__3
       (.I0(qvRAddr_WSync2[4]),
        .O(i__carry_i_1__3_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_2__3
       (.I0(qvRAddr_WSync2[3]),
        .O(i__carry_i_2__3_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_3__3
       (.I0(qvRAddr_WSync2[2]),
        .O(i__carry_i_3__3_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_4__3
       (.I0(qvRAddr_WSync2[1]),
        .O(i__carry_i_4__3_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_5__3
       (.I0(qvRAddr_WSync2[0]),
        .O(i__carry_i_5__3_n_0));
  LUT5 #(
    .INIT(32'h9A999599)) 
    i__carry_i_6__2
       (.I0(qvRAddr_WSync2[5]),
        .I1(vWAddr),
        .I2(\qvWCount_reg_n_0_[5] ),
        .I3(Q),
        .I4(qvNextWAddr_reg[5]),
        .O(i__carry_i_6__2_n_0));
  LUT5 #(
    .INIT(32'h9A999599)) 
    i__carry_i_7__2
       (.I0(qvRAddr_WSync2[4]),
        .I1(ADDRH[4]),
        .I2(\qvWCount_reg_n_0_[5] ),
        .I3(Q),
        .I4(qvNextWAddr_reg[4]),
        .O(i__carry_i_7__2_n_0));
  LUT5 #(
    .INIT(32'h9A999599)) 
    i__carry_i_8__1
       (.I0(qvRAddr_WSync2[3]),
        .I1(ADDRH[3]),
        .I2(\qvWCount_reg_n_0_[5] ),
        .I3(Q),
        .I4(qvNextWAddr_reg[3]),
        .O(i__carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h9A999599)) 
    i__carry_i_9__2
       (.I0(qvRAddr_WSync2[2]),
        .I1(ADDRH[2]),
        .I2(\qvWCount_reg_n_0_[5] ),
        .I3(Q),
        .I4(qvNextWAddr_reg[2]),
        .O(i__carry_i_9__2_n_0));
  LUT5 #(
    .INIT(32'h000F2222)) 
    qREmpty_int_i_1
       (.I0(qREmpty_int_i_2_n_0),
        .I1(qREmpty_int_i_3_n_0),
        .I2(qREmpty_int_i_4_n_0),
        .I3(qREmpty_int_i_5_n_0),
        .I4(qREmpty_int_reg_n_0),
        .O(qREmpty_int_i_1_n_0));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    qREmpty_int_i_2
       (.I0(qvPreWGrayAddr_RSync2[5]),
        .I1(qvRGrayAddr[5]),
        .I2(qvRGrayAddr[4]),
        .I3(qvPreWGrayAddr_RSync2[4]),
        .I4(qvRGrayAddr[3]),
        .I5(qvPreWGrayAddr_RSync2[3]),
        .O(qREmpty_int_i_2_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    qREmpty_int_i_3
       (.I0(qvPreWGrayAddr_RSync2[0]),
        .I1(qvRGrayAddr[0]),
        .I2(qvRGrayAddr[1]),
        .I3(qvPreWGrayAddr_RSync2[1]),
        .I4(qvRGrayAddr[2]),
        .I5(qvPreWGrayAddr_RSync2[2]),
        .O(qREmpty_int_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    qREmpty_int_i_4
       (.I0(qvRGrayAddr[5]),
        .I1(qvWGrayAddr_RSync2[5]),
        .I2(qvRGrayAddr[4]),
        .I3(qvWGrayAddr_RSync2[4]),
        .I4(qvWGrayAddr_RSync2[3]),
        .I5(qvRGrayAddr[3]),
        .O(qREmpty_int_i_4_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    qREmpty_int_i_5
       (.I0(qvWGrayAddr_RSync2[0]),
        .I1(qvRGrayAddr[0]),
        .I2(qvRGrayAddr[2]),
        .I3(qvWGrayAddr_RSync2[2]),
        .I4(qvRGrayAddr[1]),
        .I5(qvWGrayAddr_RSync2[1]),
        .O(qREmpty_int_i_5_n_0));
  FDPE #(
    .INIT(1'b1)) 
    qREmpty_int_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(qREmpty_int_i_1_n_0),
        .PRE(rst_i_0),
        .Q(qREmpty_int_reg_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    \qvDataOut[71]_i_1 
       (.I0(qREmpty_int_reg_n_0),
        .O(MemREn));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[0] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [0]),
        .Q(\qvDataOut_reg[71]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[10] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [10]),
        .Q(\qvDataOut_reg[71]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[11] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [11]),
        .Q(\qvDataOut_reg[71]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[12] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [12]),
        .Q(\qvDataOut_reg[71]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[13] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [13]),
        .Q(\qvDataOut_reg[71]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[14] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [14]),
        .Q(\qvDataOut_reg[71]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[15] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [15]),
        .Q(\qvDataOut_reg[71]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[16] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [16]),
        .Q(\qvDataOut_reg[71]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[17] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [17]),
        .Q(\qvDataOut_reg[71]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[18] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [18]),
        .Q(\qvDataOut_reg[71]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[19] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [19]),
        .Q(\qvDataOut_reg[71]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[1] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [1]),
        .Q(\qvDataOut_reg[71]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[20] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [20]),
        .Q(\qvDataOut_reg[71]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[21] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [21]),
        .Q(\qvDataOut_reg[71]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[22] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [22]),
        .Q(\qvDataOut_reg[71]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[23] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [23]),
        .Q(\qvDataOut_reg[71]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[24] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [24]),
        .Q(\qvDataOut_reg[71]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[25] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [25]),
        .Q(\qvDataOut_reg[71]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[26] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [26]),
        .Q(\qvDataOut_reg[71]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[27] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [27]),
        .Q(\qvDataOut_reg[71]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[28] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [28]),
        .Q(\qvDataOut_reg[71]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[29] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [29]),
        .Q(\qvDataOut_reg[71]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[2] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [2]),
        .Q(\qvDataOut_reg[71]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[30] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [30]),
        .Q(\qvDataOut_reg[71]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[31] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [31]),
        .Q(\qvDataOut_reg[71]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[32] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [32]),
        .Q(\qvDataOut_reg[71]_0 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[33] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [33]),
        .Q(\qvDataOut_reg[71]_0 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[34] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [34]),
        .Q(\qvDataOut_reg[71]_0 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[35] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [35]),
        .Q(\qvDataOut_reg[71]_0 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[36] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [36]),
        .Q(\qvDataOut_reg[71]_0 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[37] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [37]),
        .Q(\qvDataOut_reg[71]_0 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[38] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [38]),
        .Q(\qvDataOut_reg[71]_0 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[39] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [39]),
        .Q(\qvDataOut_reg[71]_0 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[3] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [3]),
        .Q(\qvDataOut_reg[71]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[40] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [40]),
        .Q(\qvDataOut_reg[71]_0 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[41] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [41]),
        .Q(\qvDataOut_reg[71]_0 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[42] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [42]),
        .Q(\qvDataOut_reg[71]_0 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[43] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [43]),
        .Q(\qvDataOut_reg[71]_0 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[44] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [44]),
        .Q(\qvDataOut_reg[71]_0 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[45] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [45]),
        .Q(\qvDataOut_reg[71]_0 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[46] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [46]),
        .Q(\qvDataOut_reg[71]_0 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[47] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [47]),
        .Q(\qvDataOut_reg[71]_0 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[48] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [48]),
        .Q(\qvDataOut_reg[71]_0 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[49] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [49]),
        .Q(\qvDataOut_reg[71]_0 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[4] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [4]),
        .Q(\qvDataOut_reg[71]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[50] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [50]),
        .Q(\qvDataOut_reg[71]_0 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[51] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [51]),
        .Q(\qvDataOut_reg[71]_0 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[52] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [52]),
        .Q(\qvDataOut_reg[71]_0 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[53] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [53]),
        .Q(\qvDataOut_reg[71]_0 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[54] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [54]),
        .Q(\qvDataOut_reg[71]_0 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[55] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [55]),
        .Q(\qvDataOut_reg[71]_0 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[56] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [56]),
        .Q(\qvDataOut_reg[71]_0 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[57] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [57]),
        .Q(\qvDataOut_reg[71]_0 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[58] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [58]),
        .Q(\qvDataOut_reg[71]_0 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[59] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [59]),
        .Q(\qvDataOut_reg[71]_0 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[5] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [5]),
        .Q(\qvDataOut_reg[71]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[60] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [60]),
        .Q(\qvDataOut_reg[71]_0 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[61] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [61]),
        .Q(\qvDataOut_reg[71]_0 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[62] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [62]),
        .Q(\qvDataOut_reg[71]_0 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[63] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [63]),
        .Q(\qvDataOut_reg[71]_0 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[64] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [64]),
        .Q(\qvDataOut_reg[71]_0 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[65] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [65]),
        .Q(\qvDataOut_reg[71]_0 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[66] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [66]),
        .Q(\qvDataOut_reg[71]_0 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[67] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [67]),
        .Q(\qvDataOut_reg[71]_0 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[68] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [68]),
        .Q(\qvDataOut_reg[71]_0 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[69] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [69]),
        .Q(\qvDataOut_reg[71]_0 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[6] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [6]),
        .Q(\qvDataOut_reg[71]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[70] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [70]),
        .Q(\qvDataOut_reg[71]_0 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[71] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [71]),
        .Q(\qvDataOut_reg[71]_0 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[7] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [7]),
        .Q(\qvDataOut_reg[71]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[8] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [8]),
        .Q(\qvDataOut_reg[71]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \qvDataOut_reg[9] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(\qvDataOut_reg[71]_1 [9]),
        .Q(\qvDataOut_reg[71]_0 [9]));
  LUT1 #(
    .INIT(2'h1)) 
    \qvNextRAddr[0]_i_1 
       (.I0(qvNextRAddr_reg[0]),
        .O(p_0_in__5[0]));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \qvNextRAddr[2]_i_1 
       (.I0(qvNextRAddr_reg[2]),
        .I1(qvRGrayAddr[0]),
        .I2(qvNextRAddr_reg[0]),
        .O(p_0_in__5[2]));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \qvNextRAddr[3]_i_1 
       (.I0(qvNextRAddr_reg[3]),
        .I1(qvNextRAddr_reg[0]),
        .I2(qvRGrayAddr[0]),
        .I3(qvNextRAddr_reg[2]),
        .O(p_0_in__5[3]));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \qvNextRAddr[4]_i_1 
       (.I0(qvNextRAddr_reg[4]),
        .I1(qvNextRAddr_reg[2]),
        .I2(qvRGrayAddr[0]),
        .I3(qvNextRAddr_reg[0]),
        .I4(qvNextRAddr_reg[3]),
        .O(p_0_in__5[4]));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \qvNextRAddr[5]_i_1 
       (.I0(qvNextRAddr_reg[5]),
        .I1(qvNextRAddr_reg[3]),
        .I2(qvNextRAddr_reg[0]),
        .I3(qvRGrayAddr[0]),
        .I4(qvNextRAddr_reg[2]),
        .I5(qvNextRAddr_reg[4]),
        .O(p_0_in__5[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextRAddr_reg[0] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(p_0_in__5[0]),
        .Q(qvNextRAddr_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextRAddr_reg[2] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(p_0_in__5[2]),
        .Q(qvNextRAddr_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextRAddr_reg[3] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(p_0_in__5[3]),
        .Q(qvNextRAddr_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextRAddr_reg[4] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(p_0_in__5[4]),
        .Q(qvNextRAddr_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextRAddr_reg[5] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(p_0_in__5[5]),
        .Q(qvNextRAddr_reg[5]));
  LUT1 #(
    .INIT(2'h1)) 
    \qvNextWAddr[0]_i_1 
       (.I0(qvNextWAddr_reg[0]),
        .O(p_0_in__2[0]));
  LUT2 #(
    .INIT(4'h6)) 
    \qvNextWAddr[1]_i_1 
       (.I0(qvNextWAddr_reg[0]),
        .I1(qvNextWAddr_reg[1]),
        .O(qvWGrayAddr0[0]));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \qvNextWAddr[2]_i_1 
       (.I0(qvNextWAddr_reg[2]),
        .I1(qvNextWAddr_reg[1]),
        .I2(qvNextWAddr_reg[0]),
        .O(p_0_in__2[2]));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \qvNextWAddr[3]_i_1 
       (.I0(qvNextWAddr_reg[3]),
        .I1(qvNextWAddr_reg[0]),
        .I2(qvNextWAddr_reg[1]),
        .I3(qvNextWAddr_reg[2]),
        .O(p_0_in__2[3]));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \qvNextWAddr[4]_i_1 
       (.I0(qvNextWAddr_reg[4]),
        .I1(qvNextWAddr_reg[2]),
        .I2(qvNextWAddr_reg[1]),
        .I3(qvNextWAddr_reg[0]),
        .I4(qvNextWAddr_reg[3]),
        .O(p_0_in__2[4]));
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \qvNextWAddr[5]_i_1 
       (.I0(qvNextWAddr_reg[5]),
        .I1(qvNextWAddr_reg[3]),
        .I2(qvNextWAddr_reg[0]),
        .I3(qvNextWAddr_reg[1]),
        .I4(qvNextWAddr_reg[2]),
        .I5(qvNextWAddr_reg[4]),
        .O(p_0_in__2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextWAddr_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(p_0_in__2[0]),
        .Q(qvNextWAddr_reg[0]));
  FDPE #(
    .INIT(1'b1)) 
    \qvNextWAddr_reg[1] 
       (.C(clk_i),
        .CE(E),
        .D(qvWGrayAddr0[0]),
        .PRE(rst_i_0),
        .Q(qvNextWAddr_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextWAddr_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(p_0_in__2[2]),
        .Q(qvNextWAddr_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextWAddr_reg[3] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(p_0_in__2[3]),
        .Q(qvNextWAddr_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextWAddr_reg[4] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(p_0_in__2[4]),
        .Q(qvNextWAddr_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvNextWAddr_reg[5] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(p_0_in__2[5]),
        .Q(qvNextWAddr_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(ADDRH[1]),
        .Q(qvPreWGrayAddr_RSync1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr[1]),
        .Q(qvPreWGrayAddr_RSync1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr[2]),
        .Q(qvPreWGrayAddr_RSync1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr[3]),
        .Q(qvPreWGrayAddr_RSync1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr[4]),
        .Q(qvPreWGrayAddr_RSync1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr[5]),
        .Q(qvPreWGrayAddr_RSync1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr_RSync1[0]),
        .Q(qvPreWGrayAddr_RSync2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr_RSync1[1]),
        .Q(qvPreWGrayAddr_RSync2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr_RSync1[2]),
        .Q(qvPreWGrayAddr_RSync2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr_RSync1[3]),
        .Q(qvPreWGrayAddr_RSync2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr_RSync1[4]),
        .Q(qvPreWGrayAddr_RSync2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_RSync2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvPreWGrayAddr_RSync1[5]),
        .Q(qvPreWGrayAddr_RSync2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[1]),
        .Q(qvPreWGrayAddr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[2]),
        .Q(qvPreWGrayAddr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_reg[3] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[3]),
        .Q(qvPreWGrayAddr[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_reg[4] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[4]),
        .Q(qvPreWGrayAddr[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvPreWGrayAddr_reg[5] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(vWAddr),
        .Q(qvPreWGrayAddr[5]));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \qvRAddr[0]_i_1__1 
       (.I0(qvRAddr[0]),
        .I1(qREmpty_int_reg_n_0),
        .I2(qvNextRAddr_reg[0]),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \qvRAddr[1]_i_1__1 
       (.I0(qvRAddr[1]),
        .I1(qREmpty_int_reg_n_0),
        .I2(qvRGrayAddr[0]),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \qvRAddr[2]_i_1__1 
       (.I0(qvRAddr[2]),
        .I1(qREmpty_int_reg_n_0),
        .I2(qvNextRAddr_reg[2]),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \qvRAddr[3]_i_1__1 
       (.I0(qvRAddr[3]),
        .I1(qREmpty_int_reg_n_0),
        .I2(qvNextRAddr_reg[3]),
        .O(D[3]));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \qvRAddr[4]_i_1__1 
       (.I0(qvRAddr[4]),
        .I1(qREmpty_int_reg_n_0),
        .I2(qvNextRAddr_reg[4]),
        .O(D[4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    qvRAddr_WSync20
       (.I0(qvRGrayAddr_WSync2[4]),
        .I1(qvRGrayAddr_WSync2[5]),
        .I2(qvRGrayAddr_WSync2[1]),
        .I3(qvRGrayAddr_WSync2[0]),
        .I4(qvRGrayAddr_WSync2[3]),
        .I5(qvRGrayAddr_WSync2[2]),
        .O(qvRAddr_WSync20_n_0));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \qvRAddr_WSync20_inferred__0/i_ 
       (.I0(qvRGrayAddr_WSync2[5]),
        .I1(qvRGrayAddr_WSync2[2]),
        .I2(qvRGrayAddr_WSync2[1]),
        .I3(qvRGrayAddr_WSync2[4]),
        .I4(qvRGrayAddr_WSync2[3]),
        .O(\qvRAddr_WSync20_inferred__0/i__n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \qvRAddr_WSync2[2]_i_1 
       (.I0(qvRGrayAddr_WSync2[4]),
        .I1(qvRGrayAddr_WSync2[5]),
        .I2(qvRGrayAddr_WSync2[2]),
        .I3(qvRGrayAddr_WSync2[3]),
        .O(\qvRAddr_WSync2[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \qvRAddr_WSync2[3]_i_1 
       (.I0(qvRGrayAddr_WSync2[5]),
        .I1(qvRGrayAddr_WSync2[3]),
        .I2(qvRGrayAddr_WSync2[4]),
        .O(\qvRAddr_WSync2[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRAddr_WSync2[4]_i_1 
       (.I0(qvRGrayAddr_WSync2[5]),
        .I1(qvRGrayAddr_WSync2[4]),
        .O(qvRAddr_WSync20__0));
  FDPE #(
    .INIT(1'b1)) 
    \qvRAddr_WSync2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(qvRAddr_WSync20_n_0),
        .PRE(rst_i_0),
        .Q(qvRAddr_WSync2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_WSync2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(\qvRAddr_WSync20_inferred__0/i__n_0 ),
        .Q(qvRAddr_WSync2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_WSync2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(\qvRAddr_WSync2[2]_i_1_n_0 ),
        .Q(qvRAddr_WSync2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_WSync2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(\qvRAddr_WSync2[3]_i_1_n_0 ),
        .Q(qvRAddr_WSync2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_WSync2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRAddr_WSync20__0),
        .Q(qvRAddr_WSync2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_WSync2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr_WSync2[5]),
        .Q(qvRAddr_WSync2[5]));
  FDPE #(
    .INIT(1'b1)) 
    \qvRAddr_reg[0] 
       (.C(clk_i),
        .CE(MemREn),
        .D(qvNextRAddr_reg[0]),
        .PRE(rst_i_0),
        .Q(qvRAddr[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[1] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvRGrayAddr[0]),
        .Q(qvRAddr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[2] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvNextRAddr_reg[2]),
        .Q(qvRAddr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[3] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvNextRAddr_reg[3]),
        .Q(qvRAddr[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRAddr_reg[4] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvNextRAddr_reg[4]),
        .Q(qvRAddr[4]));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRGrayAddr[0]_i_1 
       (.I0(qvNextRAddr_reg[0]),
        .I1(qvRGrayAddr[0]),
        .O(qvRGrayAddr0[0]));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRGrayAddr[1]_i_1 
       (.I0(qvRGrayAddr[0]),
        .I1(qvNextRAddr_reg[2]),
        .O(qvRGrayAddr0[1]));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRGrayAddr[2]_i_1 
       (.I0(qvNextRAddr_reg[2]),
        .I1(qvNextRAddr_reg[3]),
        .O(qvRGrayAddr0[2]));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvRGrayAddr[3]_i_1 
       (.I0(qvNextRAddr_reg[3]),
        .I1(qvNextRAddr_reg[4]),
        .O(qvRGrayAddr0[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \qvRGrayAddr[4]_i_1 
       (.I0(qvNextRAddr_reg[4]),
        .I1(qvNextRAddr_reg[5]),
        .O(qvRGrayAddr0[4]));
  FDPE #(
    .INIT(1'b1)) 
    \qvRGrayAddr_WSync1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(qvRGrayAddr[0]),
        .PRE(rst_i_0),
        .Q(qvRGrayAddr_WSync1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr[1]),
        .Q(qvRGrayAddr_WSync1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr[2]),
        .Q(qvRGrayAddr_WSync1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr[3]),
        .Q(qvRGrayAddr_WSync1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr[4]),
        .Q(qvRGrayAddr_WSync1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr[5]),
        .Q(qvRGrayAddr_WSync1[5]));
  FDPE #(
    .INIT(1'b1)) 
    \qvRGrayAddr_WSync2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(qvRGrayAddr_WSync1[0]),
        .PRE(rst_i_0),
        .Q(qvRGrayAddr_WSync2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr_WSync1[1]),
        .Q(qvRGrayAddr_WSync2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr_WSync1[2]),
        .Q(qvRGrayAddr_WSync2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr_WSync1[3]),
        .Q(qvRGrayAddr_WSync2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr_WSync1[4]),
        .Q(qvRGrayAddr_WSync2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_WSync2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvRGrayAddr_WSync1[5]),
        .Q(qvRGrayAddr_WSync2[5]));
  FDPE #(
    .INIT(1'b1)) 
    \qvRGrayAddr_reg[0] 
       (.C(clk_i),
        .CE(MemREn),
        .D(qvRGrayAddr0[0]),
        .PRE(rst_i_0),
        .Q(qvRGrayAddr[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_reg[1] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvRGrayAddr0[1]),
        .Q(qvRGrayAddr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_reg[2] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvRGrayAddr0[2]),
        .Q(qvRGrayAddr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_reg[3] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvRGrayAddr0[3]),
        .Q(qvRGrayAddr[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_reg[4] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvRGrayAddr0[4]),
        .Q(qvRGrayAddr[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvRGrayAddr_reg[5] 
       (.C(clk_i),
        .CE(MemREn),
        .CLR(rst_i_0),
        .D(qvNextRAddr_reg[5]),
        .Q(qvRGrayAddr[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \qvWAddr[4]_i_1 
       (.I0(Q),
        .I1(\qvWCount_reg_n_0_[5] ),
        .O(E));
  FDPE #(
    .INIT(1'b1)) 
    \qvWAddr_reg[0] 
       (.C(clk_i),
        .CE(E),
        .D(qvNextWAddr_reg[0]),
        .PRE(rst_i_0),
        .Q(ADDRH[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvNextWAddr_reg[1]),
        .Q(ADDRH[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvNextWAddr_reg[2]),
        .Q(ADDRH[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[3] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvNextWAddr_reg[3]),
        .Q(ADDRH[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[4] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvNextWAddr_reg[4]),
        .Q(ADDRH[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWAddr_reg[5] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvNextWAddr_reg[5]),
        .Q(vWAddr));
  FDCE #(
    .INIT(1'b0)) 
    \qvWCount_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWCount),
        .Q(\qvWCount_reg_n_0_[5] ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvWGrayAddr[1]_i_1 
       (.I0(qvNextWAddr_reg[1]),
        .I1(qvNextWAddr_reg[2]),
        .O(qvWGrayAddr0[1]));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvWGrayAddr[2]_i_1 
       (.I0(qvNextWAddr_reg[2]),
        .I1(qvNextWAddr_reg[3]),
        .O(qvWGrayAddr0[2]));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \qvWGrayAddr[3]_i_1 
       (.I0(qvNextWAddr_reg[3]),
        .I1(qvNextWAddr_reg[4]),
        .O(qvWGrayAddr0[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \qvWGrayAddr[4]_i_1 
       (.I0(qvNextWAddr_reg[4]),
        .I1(qvNextWAddr_reg[5]),
        .O(qvWGrayAddr0[4]));
  FDPE #(
    .INIT(1'b1)) 
    \qvWGrayAddr_RSync1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(qvNextWAddr_reg[1]),
        .PRE(rst_i_0),
        .Q(qvWGrayAddr_RSync1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[1]),
        .Q(qvWGrayAddr_RSync1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[2]),
        .Q(qvWGrayAddr_RSync1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[3]),
        .Q(qvWGrayAddr_RSync1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr[4]),
        .Q(qvWGrayAddr_RSync1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(vWAddr),
        .Q(qvWGrayAddr_RSync1[5]));
  FDPE #(
    .INIT(1'b1)) 
    \qvWGrayAddr_RSync2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(qvWGrayAddr_RSync1[0]),
        .PRE(rst_i_0),
        .Q(qvWGrayAddr_RSync2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr_RSync1[1]),
        .Q(qvWGrayAddr_RSync2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr_RSync1[2]),
        .Q(qvWGrayAddr_RSync2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr_RSync1[3]),
        .Q(qvWGrayAddr_RSync2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr_RSync1[4]),
        .Q(qvWGrayAddr_RSync2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_RSync2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i_0),
        .D(qvWGrayAddr_RSync1[5]),
        .Q(qvWGrayAddr_RSync2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr0[1]),
        .Q(qvWGrayAddr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr0[2]),
        .Q(qvWGrayAddr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_reg[3] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr0[3]),
        .Q(qvWGrayAddr[3]));
  FDCE #(
    .INIT(1'b0)) 
    \qvWGrayAddr_reg[4] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i_0),
        .D(qvWGrayAddr0[4]),
        .Q(qvWGrayAddr[4]));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \rxc_end_data[1]_i_1 
       (.I0(\rxc_end_data[7]_i_3_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_8_n_0 ),
        .I4(\rxc_end_data[7]_i_6_n_0 ),
        .O(\qvDataOut_reg[25]_0 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFBFB)) 
    \rxc_end_data[2]_i_1 
       (.I0(\rxc_end_data[7]_i_3_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[2]_i_2_n_0 ),
        .I4(\rxc_end_data[7]_i_8_n_0 ),
        .I5(\rxc_end_data[7]_i_6_n_0 ),
        .O(\qvDataOut_reg[25]_0 [1]));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \rxc_end_data[2]_i_2 
       (.I0(\get_e_chk[6]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [70]),
        .I2(\qvDataOut_reg[71]_0 [48]),
        .I3(\qvDataOut_reg[71]_0 [49]),
        .O(\rxc_end_data[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT5 #(
    .INIT(32'hF0F0E0F0)) 
    \rxc_end_data[4]_i_1 
       (.I0(\rxc_end_data[7]_i_5_n_0 ),
        .I1(\rxc_end_data[7]_i_3_n_0 ),
        .I2(\rxc_end_data[4]_i_2_n_0 ),
        .I3(\rxc_end_data[7]_i_4_n_0 ),
        .I4(\rxc_end_data[4]_i_3_n_0 ),
        .O(\qvDataOut_reg[25]_0 [2]));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rxc_end_data[4]_i_2 
       (.I0(\qvDataOut_reg[71]_0 [2]),
        .I1(\qvDataOut_reg[71]_0 [6]),
        .I2(\qvDataOut_reg[71]_0 [3]),
        .I3(\rxc_end_data[4]_i_4_n_0 ),
        .O(\rxc_end_data[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT5 #(
    .INIT(32'h20000000)) 
    \rxc_end_data[4]_i_3 
       (.I0(\get_e_chk[1]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [9]),
        .I2(\qvDataOut_reg[71]_0 [8]),
        .I3(\qvDataOut_reg[71]_0 [65]),
        .I4(\qvDataOut_reg[71]_0 [15]),
        .O(\rxc_end_data[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \rxc_end_data[4]_i_4 
       (.I0(\qvDataOut_reg[71]_0 [5]),
        .I1(\qvDataOut_reg[71]_0 [4]),
        .I2(\qvDataOut_reg[71]_0 [1]),
        .I3(\qvDataOut_reg[71]_0 [7]),
        .I4(\qvDataOut_reg[71]_0 [0]),
        .I5(\qvDataOut_reg[71]_0 [64]),
        .O(\rxc_end_data[4]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT4 #(
    .INIT(16'h00FB)) 
    \rxc_end_data[5]_i_1 
       (.I0(\rxc_end_data[7]_i_3_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_6_n_0 ),
        .O(\qvDataOut_reg[25]_0 [3]));
  LUT4 #(
    .INIT(16'h000B)) 
    \rxc_end_data[6]_i_1 
       (.I0(\rxc_end_data[7]_i_5_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_6_n_0 ),
        .I3(\rxc_end_data[7]_i_3_n_0 ),
        .O(\qvDataOut_reg[25]_0 [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFFFFFF)) 
    \rxc_end_data[7]_i_1 
       (.I0(\rxc_end_data[7]_i_3_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_6_n_0 ),
        .I4(\rxc_end_data[7]_i_7_n_0 ),
        .I5(\rxc_end_data[7]_i_8_n_0 ),
        .O(\qvDataOut_reg[66]_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \rxc_end_data[7]_i_10 
       (.I0(\qvDataOut_reg[71]_0 [57]),
        .I1(\qvDataOut_reg[71]_0 [62]),
        .I2(\qvDataOut_reg[71]_0 [56]),
        .I3(\qvDataOut_reg[71]_0 [63]),
        .I4(\qvDataOut_reg[71]_0 [71]),
        .I5(\get_e_chk[7]_i_2_n_0 ),
        .O(\rxc_end_data[7]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \rxc_end_data[7]_i_2 
       (.I0(\rxc_end_data[7]_i_5_n_0 ),
        .I1(\rxc_end_data[7]_i_3_n_0 ),
        .I2(\rxc_end_data[7]_i_6_n_0 ),
        .I3(\rxc_end_data[7]_i_4_n_0 ),
        .O(\qvDataOut_reg[25]_0 [5]));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \rxc_end_data[7]_i_3 
       (.I0(\qvDataOut_reg[71]_0 [66]),
        .I1(\rxc_end_data[7]_i_9_n_0 ),
        .I2(\qvDataOut_reg[71]_0 [19]),
        .I3(\qvDataOut_reg[71]_0 [18]),
        .I4(\qvDataOut_reg[71]_0 [23]),
        .I5(\qvDataOut_reg[71]_0 [16]),
        .O(\rxc_end_data[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \rxc_end_data[7]_i_4 
       (.I0(\qvDataOut_reg[71]_0 [33]),
        .I1(\qvDataOut_reg[71]_0 [38]),
        .I2(\qvDataOut_reg[71]_0 [68]),
        .I3(\qvDataOut_reg[71]_0 [32]),
        .I4(\qvDataOut_reg[71]_0 [39]),
        .I5(\get_e_chk[4]_i_2_n_0 ),
        .O(\rxc_end_data[7]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT5 #(
    .INIT(32'h20000000)) 
    \rxc_end_data[7]_i_5 
       (.I0(\get_e_chk[3]_i_2_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [25]),
        .I2(\qvDataOut_reg[71]_0 [24]),
        .I3(\qvDataOut_reg[71]_0 [26]),
        .I4(\qvDataOut_reg[71]_0 [27]),
        .O(\rxc_end_data[7]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \rxc_end_data[7]_i_6 
       (.I0(\rxc_end_data[4]_i_3_n_0 ),
        .I1(\rxc_end_data[4]_i_2_n_0 ),
        .O(\rxc_end_data[7]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT5 #(
    .INIT(32'hBAAAAAAA)) 
    \rxc_end_data[7]_i_7 
       (.I0(\rxc_end_data[7]_i_10_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [49]),
        .I2(\qvDataOut_reg[71]_0 [48]),
        .I3(\qvDataOut_reg[71]_0 [70]),
        .I4(\get_e_chk[6]_i_2_n_0 ),
        .O(\rxc_end_data[7]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rxc_end_data[7]_i_8 
       (.I0(\qvDataOut_reg[71]_0 [69]),
        .I1(\qvDataOut_reg[71]_0 [40]),
        .I2(\qvDataOut_reg[71]_0 [41]),
        .I3(\get_e_chk[5]_i_2_n_0 ),
        .O(\rxc_end_data[7]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rxc_end_data[7]_i_9 
       (.I0(\qvDataOut_reg[71]_0 [21]),
        .I1(\qvDataOut_reg[71]_0 [20]),
        .I2(\qvDataOut_reg[71]_0 [22]),
        .I3(\qvDataOut_reg[71]_0 [17]),
        .O(\rxc_end_data[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    tagged_frame_i_1
       (.I0(tagged_frame_i_2_n_0),
        .I1(tagged_frame_i_3_n_0),
        .I2(tagged_frame_i_4_n_0),
        .I3(\qvDataOut_reg[71]_0 [45]),
        .I4(\qvDataOut_reg[71]_0 [48]),
        .I5(tagged_frame_i_5_n_0),
        .O(\qvDataOut_reg[45]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    tagged_frame_i_2
       (.I0(tagged_frame_i_6_n_0),
        .I1(\qvDataOut_reg[71]_0 [35]),
        .I2(\qvDataOut_reg[71]_0 [42]),
        .I3(\qvDataOut_reg[71]_0 [47]),
        .I4(\qvDataOut_reg[71]_0 [36]),
        .I5(tagged_frame_i_7_n_0),
        .O(tagged_frame_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    tagged_frame_i_3
       (.I0(\qvDataOut_reg[71]_0 [58]),
        .I1(\qvDataOut_reg[71]_0 [57]),
        .I2(\qvDataOut_reg[71]_0 [52]),
        .I3(\qvDataOut_reg[71]_0 [59]),
        .I4(tagged_frame_i_8_n_0),
        .O(tagged_frame_i_3_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    tagged_frame_i_4
       (.I0(\qvDataOut_reg[71]_0 [38]),
        .I1(\qvDataOut_reg[71]_0 [63]),
        .I2(\qvDataOut_reg[71]_0 [33]),
        .I3(\qvDataOut_reg[71]_0 [43]),
        .O(tagged_frame_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    tagged_frame_i_5
       (.I0(\qvDataOut_reg[71]_0 [32]),
        .I1(\qvDataOut_reg[71]_0 [39]),
        .O(tagged_frame_i_5_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    tagged_frame_i_6
       (.I0(\qvDataOut_reg[71]_0 [34]),
        .I1(\qvDataOut_reg[71]_0 [51]),
        .I2(\qvDataOut_reg[71]_0 [55]),
        .I3(\qvDataOut_reg[71]_0 [61]),
        .O(tagged_frame_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    tagged_frame_i_7
       (.I0(\qvDataOut_reg[71]_0 [44]),
        .I1(\qvDataOut_reg[71]_0 [54]),
        .I2(\qvDataOut_reg[71]_0 [50]),
        .I3(\qvDataOut_reg[71]_0 [53]),
        .I4(tagged_frame_i_9_n_0),
        .O(tagged_frame_i_7_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    tagged_frame_i_8
       (.I0(\qvDataOut_reg[71]_0 [60]),
        .I1(\qvDataOut_reg[71]_0 [56]),
        .I2(\qvDataOut_reg[71]_0 [46]),
        .I3(\qvDataOut_reg[71]_0 [37]),
        .O(tagged_frame_i_8_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    tagged_frame_i_9
       (.I0(\qvDataOut_reg[71]_0 [41]),
        .I1(\qvDataOut_reg[71]_0 [40]),
        .I2(\qvDataOut_reg[71]_0 [49]),
        .I3(\qvDataOut_reg[71]_0 [62]),
        .O(tagged_frame_i_9_n_0));
  LUT6 #(
    .INIT(64'hFFFF00F400000000)) 
    \terminator_location[0]_i_1 
       (.I0(\terminator_location[0]_i_2_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_3_n_0 ),
        .I4(\rxc_end_data[4]_i_3_n_0 ),
        .I5(\rxc_end_data[4]_i_2_n_0 ),
        .O(\qvDataOut_reg[69]_0 [0]));
  LUT3 #(
    .INIT(8'h8A)) 
    \terminator_location[0]_i_2 
       (.I0(\rxc_end_data[7]_i_8_n_0 ),
        .I1(\terminator_location[0]_i_3_n_0 ),
        .I2(\rxc_end_data[7]_i_10_n_0 ),
        .O(\terminator_location[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \terminator_location[0]_i_3 
       (.I0(\qvDataOut_reg[71]_0 [49]),
        .I1(\qvDataOut_reg[71]_0 [54]),
        .I2(\qvDataOut_reg[71]_0 [50]),
        .I3(\qvDataOut_reg[71]_0 [51]),
        .I4(\terminator_location[0]_i_4_n_0 ),
        .O(\terminator_location[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \terminator_location[0]_i_4 
       (.I0(\qvDataOut_reg[71]_0 [53]),
        .I1(\qvDataOut_reg[71]_0 [52]),
        .I2(\qvDataOut_reg[71]_0 [55]),
        .I3(\qvDataOut_reg[71]_0 [70]),
        .I4(\qvDataOut_reg[71]_0 [48]),
        .O(\terminator_location[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF8F0)) 
    \terminator_location[1]_i_1 
       (.I0(\rxc_end_data[7]_i_7_n_0 ),
        .I1(\terminator_location[1]_i_2_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_4_n_0 ),
        .I4(\rxc_end_data[7]_i_3_n_0 ),
        .I5(\rxc_end_data[7]_i_6_n_0 ),
        .O(\qvDataOut_reg[69]_0 [1]));
  LUT5 #(
    .INIT(32'hEFFFFFFF)) 
    \terminator_location[1]_i_2 
       (.I0(\terminator_location[1]_i_3_n_0 ),
        .I1(\qvDataOut_reg[71]_0 [41]),
        .I2(\qvDataOut_reg[71]_0 [46]),
        .I3(\qvDataOut_reg[71]_0 [42]),
        .I4(\qvDataOut_reg[71]_0 [43]),
        .O(\terminator_location[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \terminator_location[1]_i_3 
       (.I0(\qvDataOut_reg[71]_0 [45]),
        .I1(\qvDataOut_reg[71]_0 [44]),
        .I2(\qvDataOut_reg[71]_0 [47]),
        .I3(\qvDataOut_reg[71]_0 [69]),
        .I4(\qvDataOut_reg[71]_0 [40]),
        .O(\terminator_location[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000D0F)) 
    \terminator_location[2]_i_1 
       (.I0(\rxc_end_data[7]_i_8_n_0 ),
        .I1(\rxc_end_data[7]_i_7_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_4_n_0 ),
        .I4(\rxc_end_data[7]_i_3_n_0 ),
        .I5(\rxc_end_data[7]_i_6_n_0 ),
        .O(\qvDataOut_reg[69]_0 [2]));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    this_cycle_i_1
       (.I0(\rxc_end_data[7]_i_3_n_0 ),
        .I1(\rxc_end_data[7]_i_4_n_0 ),
        .I2(\rxc_end_data[7]_i_5_n_0 ),
        .I3(\rxc_end_data[7]_i_6_n_0 ),
        .O(this_cycle));
endmodule

(* ORIG_REF_NAME = "LPF3x8" *) 
module switch_elements_LPF3x8
   (d4_30,
    DO,
    clk_i,
    rst_i,
    \d4_4_reg[15]_0 ,
    FREQ,
    DI,
    E,
    out);
  output d4_30;
  output [15:0]DO;
  input clk_i;
  input rst_i;
  input \d4_4_reg[15]_0 ;
  input [11:0]FREQ;
  input [15:0]DI;
  input [0:0]E;
  input out;

  wire [17:0]A;
  wire [15:0]D;
  wire [15:0]DI;
  wire [15:0]DO;
  wire \DO[15]_i_1_n_0 ;
  wire DZ1_n_16;
  wire DZ1_n_17;
  wire DZ1_n_18;
  wire DZ1_n_19;
  wire DZ1_n_20;
  wire DZ1_n_21;
  wire DZ1_n_22;
  wire DZ1_n_23;
  wire DZ1_n_24;
  wire DZ1_n_25;
  wire DZ1_n_26;
  wire DZ1_n_27;
  wire DZ1_n_28;
  wire DZ1_n_29;
  wire DZ1_n_30;
  wire DZ1_n_31;
  wire DZ1_n_32;
  wire DZ1_n_33;
  wire DZ2_78_n_0;
  wire DZ2_78_n_1;
  wire DZ2_78_n_10;
  wire DZ2_78_n_11;
  wire DZ2_78_n_12;
  wire DZ2_78_n_13;
  wire DZ2_78_n_14;
  wire DZ2_78_n_15;
  wire DZ2_78_n_2;
  wire DZ2_78_n_3;
  wire DZ2_78_n_4;
  wire DZ2_78_n_5;
  wire DZ2_78_n_6;
  wire DZ2_78_n_7;
  wire DZ2_78_n_8;
  wire DZ2_78_n_9;
  wire DZ3_78_n_1;
  wire DZ3_78_n_10;
  wire DZ3_78_n_11;
  wire DZ3_78_n_12;
  wire DZ3_78_n_13;
  wire DZ3_78_n_14;
  wire DZ3_78_n_15;
  wire DZ3_78_n_16;
  wire DZ3_78_n_2;
  wire DZ3_78_n_3;
  wire DZ3_78_n_4;
  wire DZ3_78_n_5;
  wire DZ3_78_n_6;
  wire DZ3_78_n_7;
  wire DZ3_78_n_8;
  wire DZ3_78_n_9;
  wire DZ3_n_16;
  wire DZ3_n_17;
  wire DZ3_n_18;
  wire DZ3_n_19;
  wire DZ3_n_20;
  wire DZ3_n_21;
  wire DZ3_n_22;
  wire DZ3_n_23;
  wire DZ3_n_24;
  wire DZ3_n_25;
  wire DZ3_n_26;
  wire DZ3_n_27;
  wire DZ3_n_28;
  wire DZ3_n_29;
  wire DZ3_n_30;
  wire DZ3_n_31;
  wire DZ3_n_32;
  wire DZ3_n_33;
  wire DZ4_56_n_0;
  wire DZ4_56_n_1;
  wire DZ4_56_n_10;
  wire DZ4_56_n_11;
  wire DZ4_56_n_12;
  wire DZ4_56_n_13;
  wire DZ4_56_n_14;
  wire DZ4_56_n_15;
  wire DZ4_56_n_2;
  wire DZ4_56_n_3;
  wire DZ4_56_n_4;
  wire DZ4_56_n_5;
  wire DZ4_56_n_6;
  wire DZ4_56_n_7;
  wire DZ4_56_n_8;
  wire DZ4_56_n_9;
  wire DZ4_n_18;
  wire [0:0]E;
  wire [11:0]FREQ;
  wire [27:9]L;
  wire [15:0]Q;
  wire [19:0]R;
  wire SE;
  wire SE11_out;
  wire U_C_n_40;
  wire [11:0]a0;
  wire [11:0]a0d;
  wire [11:0]a1;
  wire a14;
  wire [11:0]a1d;
  wire activity_blocks_gate__72_n_0;
  wire activity_blocks_gate__73_n_0;
  wire activity_blocks_gate__74_n_0;
  wire activity_blocks_gate__75_n_0;
  wire activity_blocks_gate__76_n_0;
  wire activity_blocks_gate__77_n_0;
  wire activity_blocks_gate__78_n_0;
  wire activity_blocks_gate__79_n_0;
  wire activity_blocks_gate__80_n_0;
  wire activity_blocks_gate__81_n_0;
  wire activity_blocks_gate__82_n_0;
  wire activity_blocks_gate__83_n_0;
  wire activity_blocks_gate__84_n_0;
  wire activity_blocks_gate__85_n_0;
  wire activity_blocks_gate__86_n_0;
  wire activity_blocks_gate__87_n_0;
  wire [11:0]b1;
  wire [11:0]b1d;
  wire clk_i;
  wire [15:0]d1_3;
  wire [15:0]d1_4;
  wire [15:0]d2_3;
  wire [15:0]d2_4;
  wire [15:0]d3_3;
  wire [15:0]d3_4;
  wire d4_30;
  wire \d4_3_reg[0]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[10]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[11]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[12]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[13]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[14]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[15]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[1]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[2]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[3]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[4]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[5]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[6]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[7]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[8]_srl2_activity_blocks_c_10_n_0 ;
  wire \d4_3_reg[9]_srl2_activity_blocks_c_10_n_0 ;
  wire [15:0]d4_4;
  wire \d4_40_reg[0]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[10]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[11]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[12]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[13]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[14]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[15]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[1]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[2]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[3]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[4]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[5]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[6]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[7]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[8]_activity_blocks_c_11_n_0 ;
  wire \d4_40_reg[9]_activity_blocks_c_11_n_0 ;
  wire \d4_4_reg[15]_0 ;
  wire [15:0]d56_2;
  wire [15:0]d56_3;
  wire [15:0]d78_1;
  wire [15:0]d78_2;
  wire [15:0]d78_3;
  wire \d_z2[20]_i_2_n_0 ;
  wire \d_z2[20]_i_3_n_0 ;
  wire \d_z2[20]_i_4_n_0 ;
  wire \d_z2[20]_i_5_n_0 ;
  wire \d_z2[20]_i_6_n_0 ;
  wire [18:0]dd1;
  wire [15:0]dd2;
  wire [18:16]dd2__0;
  wire [15:0]did;
  wire \did[15]_i_1_n_0 ;
  wire [18:0]dii;
  wire doii1;
  wire [20:3]minusOp;
  wire out;
  wire [15:14]p_1_in__0;
  wire [18:0]plusOp;
  wire [18:17]plusOp18;
  wire rst_i;
  wire [0:0]sh;
  wire [2:0]st;
  wire \st[0]_i_1__0_n_0 ;
  wire \st[1]_i_1__0_n_0 ;
  wire \st[2]_i_1__0_n_0 ;
  wire t1_reg_n_100;
  wire t1_reg_n_101;
  wire t1_reg_n_102;
  wire t1_reg_n_103;
  wire t1_reg_n_104;
  wire t1_reg_n_105;
  wire t1_reg_n_77;
  wire t1_reg_n_78;
  wire t1_reg_n_79;
  wire t1_reg_n_80;
  wire t1_reg_n_81;
  wire t1_reg_n_82;
  wire t1_reg_n_83;
  wire t1_reg_n_84;
  wire t1_reg_n_85;
  wire t1_reg_n_86;
  wire t1_reg_n_87;
  wire t1_reg_n_88;
  wire t1_reg_n_89;
  wire t1_reg_n_90;
  wire t1_reg_n_91;
  wire t1_reg_n_92;
  wire t1_reg_n_93;
  wire t1_reg_n_94;
  wire t1_reg_n_95;
  wire t1_reg_n_96;
  wire t1_reg_n_97;
  wire t1_reg_n_98;
  wire t1_reg_n_99;
  wire t2_reg_n_100;
  wire t2_reg_n_101;
  wire t2_reg_n_102;
  wire t2_reg_n_103;
  wire t2_reg_n_104;
  wire t2_reg_n_105;
  wire t2_reg_n_77;
  wire t2_reg_n_98;
  wire t2_reg_n_99;
  wire [19:0]t2z2;
  wire \t2z2[15]_i_2_n_0 ;
  wire \t2z2[15]_i_3_n_0 ;
  wire \t2z2[15]_i_4_n_0 ;
  wire \t2z2[15]_i_5_n_0 ;
  wire \t2z2[15]_i_6_n_0 ;
  wire \t2z2[15]_i_7_n_0 ;
  wire \t2z2[15]_i_8_n_0 ;
  wire \t2z2[15]_i_9_n_0 ;
  wire \t2z2[7]_i_2_n_0 ;
  wire \t2z2[7]_i_3_n_0 ;
  wire \t2z2[7]_i_4_n_0 ;
  wire \t2z2[7]_i_5_n_0 ;
  wire \t2z2[7]_i_6_n_0 ;
  wire \t2z2[7]_i_7_n_0 ;
  wire \t2z2[7]_i_8_n_0 ;
  wire \t2z2[7]_i_9_n_0 ;
  wire \t2z2_reg[15]_i_1_n_0 ;
  wire \t2z2_reg[15]_i_1_n_1 ;
  wire \t2z2_reg[15]_i_1_n_2 ;
  wire \t2z2_reg[15]_i_1_n_3 ;
  wire \t2z2_reg[15]_i_1_n_4 ;
  wire \t2z2_reg[15]_i_1_n_5 ;
  wire \t2z2_reg[15]_i_1_n_6 ;
  wire \t2z2_reg[15]_i_1_n_7 ;
  wire \t2z2_reg[19]_i_1_n_5 ;
  wire \t2z2_reg[19]_i_1_n_6 ;
  wire \t2z2_reg[19]_i_1_n_7 ;
  wire \t2z2_reg[7]_i_1_n_0 ;
  wire \t2z2_reg[7]_i_1_n_1 ;
  wire \t2z2_reg[7]_i_1_n_2 ;
  wire \t2z2_reg[7]_i_1_n_3 ;
  wire \t2z2_reg[7]_i_1_n_4 ;
  wire \t2z2_reg[7]_i_1_n_5 ;
  wire \t2z2_reg[7]_i_1_n_6 ;
  wire \t2z2_reg[7]_i_1_n_7 ;
  wire [19:2]t2z2_z3;
  wire \t2z2_z3[19]_i_2_n_0 ;
  wire \t2z2_z3[19]_i_3_n_0 ;
  wire \t2z2_z3[19]_i_4_n_0 ;
  wire \t2z2_z3[19]_i_5_n_0 ;
  wire [15:0]t2z2d1;
  wire [15:0]t2z2d2;
  wire [19:0]t2z2i;
  wire t3_reg_n_100;
  wire t3_reg_n_101;
  wire t3_reg_n_102;
  wire t3_reg_n_103;
  wire t3_reg_n_104;
  wire t3_reg_n_105;
  wire t3_reg_n_77;
  wire t3_reg_n_97;
  wire t3_reg_n_98;
  wire t3_reg_n_99;
  wire [18:0]t3z3;
  wire \t3z3[15]_i_2_n_0 ;
  wire \t3z3[15]_i_3_n_0 ;
  wire \t3z3[15]_i_4_n_0 ;
  wire \t3z3[15]_i_5_n_0 ;
  wire \t3z3[15]_i_6_n_0 ;
  wire \t3z3[15]_i_7_n_0 ;
  wire \t3z3[15]_i_8_n_0 ;
  wire \t3z3[15]_i_9_n_0 ;
  wire \t3z3[7]_i_2_n_0 ;
  wire \t3z3[7]_i_3_n_0 ;
  wire \t3z3[7]_i_4_n_0 ;
  wire \t3z3[7]_i_5_n_0 ;
  wire \t3z3[7]_i_6_n_0 ;
  wire \t3z3[7]_i_7_n_0 ;
  wire \t3z3[7]_i_8_n_0 ;
  wire \t3z3[7]_i_9_n_0 ;
  wire \t3z3_reg[15]_i_1_n_0 ;
  wire \t3z3_reg[15]_i_1_n_1 ;
  wire \t3z3_reg[15]_i_1_n_2 ;
  wire \t3z3_reg[15]_i_1_n_3 ;
  wire \t3z3_reg[15]_i_1_n_4 ;
  wire \t3z3_reg[15]_i_1_n_5 ;
  wire \t3z3_reg[15]_i_1_n_6 ;
  wire \t3z3_reg[15]_i_1_n_7 ;
  wire \t3z3_reg[18]_i_1_n_6 ;
  wire \t3z3_reg[18]_i_1_n_7 ;
  wire \t3z3_reg[7]_i_1_n_0 ;
  wire \t3z3_reg[7]_i_1_n_1 ;
  wire \t3z3_reg[7]_i_1_n_2 ;
  wire \t3z3_reg[7]_i_1_n_3 ;
  wire \t3z3_reg[7]_i_1_n_4 ;
  wire \t3z3_reg[7]_i_1_n_5 ;
  wire \t3z3_reg[7]_i_1_n_6 ;
  wire \t3z3_reg[7]_i_1_n_7 ;
  wire [15:0]tt1;
  wire [20:0]tt2;
  wire \tt2[15]_i_2_n_0 ;
  wire \tt2[15]_i_3_n_0 ;
  wire \tt2[15]_i_4_n_0 ;
  wire \tt2[15]_i_5_n_0 ;
  wire \tt2[15]_i_6_n_0 ;
  wire \tt2[15]_i_7_n_0 ;
  wire \tt2[15]_i_8_n_0 ;
  wire \tt2[15]_i_9_n_0 ;
  wire \tt2[20]_i_2_n_0 ;
  wire \tt2[20]_i_3_n_0 ;
  wire \tt2[20]_i_4_n_0 ;
  wire \tt2[20]_i_5_n_0 ;
  wire \tt2[20]_i_6_n_0 ;
  wire \tt2[20]_i_7_n_0 ;
  wire \tt2[7]_i_2_n_0 ;
  wire \tt2[7]_i_3_n_0 ;
  wire \tt2[7]_i_4_n_0 ;
  wire \tt2[7]_i_5_n_0 ;
  wire \tt2[7]_i_6_n_0 ;
  wire \tt2[7]_i_7_n_0 ;
  wire \tt2[7]_i_8_n_0 ;
  wire \tt2[7]_i_9_n_0 ;
  wire \tt2_reg[15]_i_1_n_0 ;
  wire \tt2_reg[15]_i_1_n_1 ;
  wire \tt2_reg[15]_i_1_n_10 ;
  wire \tt2_reg[15]_i_1_n_11 ;
  wire \tt2_reg[15]_i_1_n_12 ;
  wire \tt2_reg[15]_i_1_n_13 ;
  wire \tt2_reg[15]_i_1_n_14 ;
  wire \tt2_reg[15]_i_1_n_15 ;
  wire \tt2_reg[15]_i_1_n_2 ;
  wire \tt2_reg[15]_i_1_n_3 ;
  wire \tt2_reg[15]_i_1_n_4 ;
  wire \tt2_reg[15]_i_1_n_5 ;
  wire \tt2_reg[15]_i_1_n_6 ;
  wire \tt2_reg[15]_i_1_n_7 ;
  wire \tt2_reg[15]_i_1_n_8 ;
  wire \tt2_reg[15]_i_1_n_9 ;
  wire \tt2_reg[20]_i_1_n_11 ;
  wire \tt2_reg[20]_i_1_n_12 ;
  wire \tt2_reg[20]_i_1_n_13 ;
  wire \tt2_reg[20]_i_1_n_14 ;
  wire \tt2_reg[20]_i_1_n_15 ;
  wire \tt2_reg[20]_i_1_n_4 ;
  wire \tt2_reg[20]_i_1_n_5 ;
  wire \tt2_reg[20]_i_1_n_6 ;
  wire \tt2_reg[20]_i_1_n_7 ;
  wire \tt2_reg[7]_i_1_n_0 ;
  wire \tt2_reg[7]_i_1_n_1 ;
  wire \tt2_reg[7]_i_1_n_10 ;
  wire \tt2_reg[7]_i_1_n_11 ;
  wire \tt2_reg[7]_i_1_n_12 ;
  wire \tt2_reg[7]_i_1_n_13 ;
  wire \tt2_reg[7]_i_1_n_14 ;
  wire \tt2_reg[7]_i_1_n_15 ;
  wire \tt2_reg[7]_i_1_n_2 ;
  wire \tt2_reg[7]_i_1_n_3 ;
  wire \tt2_reg[7]_i_1_n_4 ;
  wire \tt2_reg[7]_i_1_n_5 ;
  wire \tt2_reg[7]_i_1_n_6 ;
  wire \tt2_reg[7]_i_1_n_7 ;
  wire \tt2_reg[7]_i_1_n_8 ;
  wire \tt2_reg[7]_i_1_n_9 ;
  wire [21:4]tt2_z1;
  wire \tt2_z1[21]_i_2_n_0 ;
  wire \tt2_z1[21]_i_3_n_0 ;
  wire \tt2_z1[21]_i_4_n_0 ;
  wire \tt2_z1[21]_i_5_n_0 ;
  wire \tt2_z1[21]_i_6_n_0 ;
  wire [15:0]tt2d1;
  wire [15:0]tt2d2;
  wire [15:0]z1;
  wire [15:0]z1d1;
  wire [15:0]z1d2;
  wire [15:0]z1i;
  wire [15:0]z2;
  wire [15:0]z2d1;
  wire [15:0]z2d2;
  wire [15:0]z2i;
  wire [15:0]z3;
  wire [15:0]z3d1;
  wire [15:0]z3d2;
  wire [15:0]z3i;
  wire [15:0]z4i;
  wire NLW_t1_reg_CARRYCASCOUT_UNCONNECTED;
  wire NLW_t1_reg_MULTSIGNOUT_UNCONNECTED;
  wire NLW_t1_reg_OVERFLOW_UNCONNECTED;
  wire NLW_t1_reg_PATTERNBDETECT_UNCONNECTED;
  wire NLW_t1_reg_PATTERNDETECT_UNCONNECTED;
  wire NLW_t1_reg_UNDERFLOW_UNCONNECTED;
  wire [29:0]NLW_t1_reg_ACOUT_UNCONNECTED;
  wire [17:0]NLW_t1_reg_BCOUT_UNCONNECTED;
  wire [3:0]NLW_t1_reg_CARRYOUT_UNCONNECTED;
  wire [47:29]NLW_t1_reg_P_UNCONNECTED;
  wire [47:0]NLW_t1_reg_PCOUT_UNCONNECTED;
  wire [7:0]NLW_t1_reg_XOROUT_UNCONNECTED;
  wire NLW_t2_reg_CARRYCASCOUT_UNCONNECTED;
  wire NLW_t2_reg_MULTSIGNOUT_UNCONNECTED;
  wire NLW_t2_reg_OVERFLOW_UNCONNECTED;
  wire NLW_t2_reg_PATTERNBDETECT_UNCONNECTED;
  wire NLW_t2_reg_PATTERNDETECT_UNCONNECTED;
  wire NLW_t2_reg_UNDERFLOW_UNCONNECTED;
  wire [29:0]NLW_t2_reg_ACOUT_UNCONNECTED;
  wire [17:0]NLW_t2_reg_BCOUT_UNCONNECTED;
  wire [3:0]NLW_t2_reg_CARRYOUT_UNCONNECTED;
  wire [47:29]NLW_t2_reg_P_UNCONNECTED;
  wire [47:0]NLW_t2_reg_PCOUT_UNCONNECTED;
  wire [7:0]NLW_t2_reg_XOROUT_UNCONNECTED;
  wire [7:3]\NLW_t2z2_reg[19]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_t2z2_reg[19]_i_1_O_UNCONNECTED ;
  wire NLW_t3_reg_CARRYCASCOUT_UNCONNECTED;
  wire NLW_t3_reg_MULTSIGNOUT_UNCONNECTED;
  wire NLW_t3_reg_OVERFLOW_UNCONNECTED;
  wire NLW_t3_reg_PATTERNBDETECT_UNCONNECTED;
  wire NLW_t3_reg_PATTERNDETECT_UNCONNECTED;
  wire NLW_t3_reg_UNDERFLOW_UNCONNECTED;
  wire [29:0]NLW_t3_reg_ACOUT_UNCONNECTED;
  wire [17:0]NLW_t3_reg_BCOUT_UNCONNECTED;
  wire [3:0]NLW_t3_reg_CARRYOUT_UNCONNECTED;
  wire [47:29]NLW_t3_reg_P_UNCONNECTED;
  wire [47:0]NLW_t3_reg_PCOUT_UNCONNECTED;
  wire [7:0]NLW_t3_reg_XOROUT_UNCONNECTED;
  wire [7:2]\NLW_t3z3_reg[18]_i_1_CO_UNCONNECTED ;
  wire [7:3]\NLW_t3z3_reg[18]_i_1_O_UNCONNECTED ;
  wire [7:4]\NLW_tt2_reg[20]_i_1_CO_UNCONNECTED ;
  wire [7:5]\NLW_tt2_reg[20]_i_1_O_UNCONNECTED ;

  switch_elements_DELAY__parameterized20 DD
       (.D(dii[15:0]),
        .DI({\d_z2[20]_i_2_n_0 ,\d_z2[20]_i_3_n_0 }),
        .Q(st),
        .S({\d_z2[20]_i_4_n_0 ,\d_z2[20]_i_5_n_0 ,\d_z2[20]_i_6_n_0 }),
        .clk_i(clk_i),
        .\d_z2_reg[15] (z2),
        .\dd1_reg[15] (did[13:0]),
        .\dd1_reg[15]_0 (D),
        .\did_reg[15] ({minusOp[20],minusOp[18:3]}));
  LUT3 #(
    .INIT(8'h08)) 
    \DO[15]_i_1 
       (.I0(st[2]),
        .I1(st[1]),
        .I2(st[0]),
        .O(\DO[15]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[0] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[2]),
        .Q(DO[0]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[10] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[12]),
        .Q(DO[10]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[11] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[13]),
        .Q(DO[11]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[12] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[14]),
        .Q(DO[12]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[13] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[15]),
        .Q(DO[13]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[14] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_1_in__0[14]),
        .Q(DO[14]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[15] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_1_in__0[15]),
        .Q(DO[15]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[1] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[3]),
        .Q(DO[1]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[2] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[4]),
        .Q(DO[2]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[3] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[5]),
        .Q(DO[3]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[4] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[6]),
        .Q(DO[4]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[5] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[7]),
        .Q(DO[5]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[6] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[8]),
        .Q(DO[6]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[7] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[9]),
        .Q(DO[7]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[8] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[10]),
        .Q(DO[8]));
  FDCE #(
    .INIT(1'b0)) 
    \DO_reg[9] 
       (.C(clk_i),
        .CE(\DO[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(D[11]),
        .Q(DO[9]));
  switch_elements_DELAY DZ1
       (.D({DZ1_n_16,DZ1_n_17,DZ1_n_18,DZ1_n_19,DZ1_n_20,DZ1_n_21,DZ1_n_22,DZ1_n_23,DZ1_n_24,DZ1_n_25,DZ1_n_26,DZ1_n_27,DZ1_n_28,DZ1_n_29,DZ1_n_30,DZ1_n_31,DZ1_n_32,DZ1_n_33}),
        .Q(tt2[19:0]),
        .S({\tt2_z1[21]_i_2_n_0 ,\tt2_z1[21]_i_3_n_0 ,\tt2_z1[21]_i_4_n_0 ,\tt2_z1[21]_i_5_n_0 ,\tt2_z1[21]_i_6_n_0 }),
        .clk_i(clk_i),
        .clk_i_0(z1),
        .\z1d1_reg[15] (z1i));
  switch_elements_DELAY_0 DZ1_56
       (.D(tt1),
        .Q(Q),
        .SE11_out(SE11_out),
        .clk_i(clk_i));
  switch_elements_DELAY__parameterized7 DZ1_78
       (.D(tt1),
        .P({t1_reg_n_83,t1_reg_n_84,t1_reg_n_85,t1_reg_n_86,t1_reg_n_87,t1_reg_n_88,t1_reg_n_89,t1_reg_n_90,t1_reg_n_91,t1_reg_n_92,t1_reg_n_93,t1_reg_n_94,t1_reg_n_95,t1_reg_n_96,t1_reg_n_97,t1_reg_n_98}),
        .Q(tt2d2),
        .SE(SE),
        .clk_i(clk_i),
        .clk_i_0(d78_1));
  switch_elements_DELAY__parameterized16 DZ2
       (.D(z2i),
        .Q(z2),
        .clk_i(clk_i));
  switch_elements_DELAY__parameterized1 DZ2_56
       (.D({DZ2_78_n_0,DZ2_78_n_1,DZ2_78_n_2,DZ2_78_n_3,DZ2_78_n_4,DZ2_78_n_5,DZ2_78_n_6,DZ2_78_n_7,DZ2_78_n_8,DZ2_78_n_9,DZ2_78_n_10,DZ2_78_n_11,DZ2_78_n_12,DZ2_78_n_13,DZ2_78_n_14,DZ2_78_n_15}),
        .Q(d56_2),
        .SE11_out(SE11_out),
        .clk_i(clk_i));
  switch_elements_DELAY__parameterized9 DZ2_78
       (.D({DZ2_78_n_0,DZ2_78_n_1,DZ2_78_n_2,DZ2_78_n_3,DZ2_78_n_4,DZ2_78_n_5,DZ2_78_n_6,DZ2_78_n_7,DZ2_78_n_8,DZ2_78_n_9,DZ2_78_n_10,DZ2_78_n_11,DZ2_78_n_12,DZ2_78_n_13,DZ2_78_n_14,DZ2_78_n_15}),
        .P({t1_reg_n_83,t1_reg_n_84,t1_reg_n_85,t1_reg_n_86,t1_reg_n_87,t1_reg_n_88,t1_reg_n_89,t1_reg_n_90,t1_reg_n_91,t1_reg_n_92,t1_reg_n_93,t1_reg_n_94,t1_reg_n_95,t1_reg_n_96,t1_reg_n_97,t1_reg_n_98}),
        .Q(z1d2),
        .SE(SE),
        .clk_i(clk_i),
        .clk_i_0(d78_2));
  switch_elements_DELAY__parameterized3 DZ3
       (.D({DZ3_n_16,DZ3_n_17,DZ3_n_18,DZ3_n_19,DZ3_n_20,DZ3_n_21,DZ3_n_22,DZ3_n_23,DZ3_n_24,DZ3_n_25,DZ3_n_26,DZ3_n_27,DZ3_n_28,DZ3_n_29,DZ3_n_30,DZ3_n_31,DZ3_n_32,DZ3_n_33}),
        .Q(t2z2[18:0]),
        .S({\t2z2_z3[19]_i_2_n_0 ,\t2z2_z3[19]_i_3_n_0 ,\t2z2_z3[19]_i_4_n_0 ,\t2z2_z3[19]_i_5_n_0 }),
        .clk_i(clk_i),
        .clk_i_0(z3),
        .\z3d1_reg[15] (z3i));
  switch_elements_DELAY__parameterized3_1 DZ3_56
       (.D({DZ3_78_n_1,DZ3_78_n_2,DZ3_78_n_3,DZ3_78_n_4,DZ3_78_n_5,DZ3_78_n_6,DZ3_78_n_7,DZ3_78_n_8,DZ3_78_n_9,DZ3_78_n_10,DZ3_78_n_11,DZ3_78_n_12,DZ3_78_n_13,DZ3_78_n_14,DZ3_78_n_15,DZ3_78_n_16}),
        .Q(st[2:1]),
        .SE11_out(SE11_out),
        .clk_i(clk_i),
        .clk_i_0(d56_3));
  switch_elements_DELAY__parameterized11 DZ3_78
       (.D({DZ3_78_n_1,DZ3_78_n_2,DZ3_78_n_3,DZ3_78_n_4,DZ3_78_n_5,DZ3_78_n_6,DZ3_78_n_7,DZ3_78_n_8,DZ3_78_n_9,DZ3_78_n_10,DZ3_78_n_11,DZ3_78_n_12,DZ3_78_n_13,DZ3_78_n_14,DZ3_78_n_15,DZ3_78_n_16}),
        .P(L[24:9]),
        .Q(st[2:1]),
        .SE(SE),
        .clk_i(clk_i),
        .clk_i_0(d78_3),
        .\d3_3_reg[15] (t2z2d2));
  switch_elements_DELAY__parameterized18 DZ4
       (.D(z4i),
        .\DO_reg[15] (t3z3),
        .O(plusOp18),
        .Q(st),
        .clk_i(clk_i),
        .clk_i_0(D),
        .doii1(doii1),
        .\st_reg[2] (DZ4_n_18));
  switch_elements_DELAY__parameterized5 DZ4_56
       (.\D32.DEL1[15].U_SRL0_i_1 (dd2),
        .\D32.DEL1[15].U_SRL0_i_1_0 (sh),
        .Q(st),
        .clk_i(clk_i),
        .\dd2_reg[0] (DZ4_56_n_0),
        .\dd2_reg[10] (DZ4_56_n_10),
        .\dd2_reg[11] (DZ4_56_n_11),
        .\dd2_reg[12] (DZ4_56_n_12),
        .\dd2_reg[13] (DZ4_56_n_13),
        .\dd2_reg[14] (DZ4_56_n_14),
        .\dd2_reg[15] (DZ4_56_n_15),
        .\dd2_reg[1] (DZ4_56_n_1),
        .\dd2_reg[2] (DZ4_56_n_2),
        .\dd2_reg[3] (DZ4_56_n_3),
        .\dd2_reg[4] (DZ4_56_n_4),
        .\dd2_reg[5] (DZ4_56_n_5),
        .\dd2_reg[6] (DZ4_56_n_6),
        .\dd2_reg[7] (DZ4_56_n_7),
        .\dd2_reg[8] (DZ4_56_n_8),
        .\dd2_reg[9] (DZ4_56_n_9));
  switch_elements_DELAY__parameterized13 DZ4_78
       (.D(z4i),
        .\D32.DEL1[0].U_SRL0_0 (DZ4_56_n_0),
        .\D32.DEL1[10].U_SRL0_0 (DZ4_56_n_10),
        .\D32.DEL1[11].U_SRL0_0 (DZ4_56_n_11),
        .\D32.DEL1[12].U_SRL0_0 (DZ4_56_n_12),
        .\D32.DEL1[13].U_SRL0_0 (DZ4_56_n_13),
        .\D32.DEL1[14].U_SRL0_0 (DZ4_56_n_14),
        .\D32.DEL1[15].U_SRL0_0 (DZ4_n_18),
        .\D32.DEL1[15].U_SRL0_1 (U_C_n_40),
        .\D32.DEL1[15].U_SRL0_2 (DZ4_56_n_15),
        .\D32.DEL1[15].U_SRL1_0 (dd2),
        .\D32.DEL1[1].U_SRL0_0 (DZ4_56_n_1),
        .\D32.DEL1[2].U_SRL0_0 (DZ4_56_n_2),
        .\D32.DEL1[3].U_SRL0_0 (DZ4_56_n_3),
        .\D32.DEL1[4].U_SRL0_0 (DZ4_56_n_4),
        .\D32.DEL1[5].U_SRL0_0 (DZ4_56_n_5),
        .\D32.DEL1[6].U_SRL0_0 (DZ4_56_n_6),
        .\D32.DEL1[7].U_SRL0_0 (DZ4_56_n_7),
        .\D32.DEL1[8].U_SRL0_0 (DZ4_56_n_8),
        .\D32.DEL1[9].U_SRL0_0 (DZ4_56_n_9),
        .Q(st),
        .clk_i(clk_i),
        .d4_4(d4_4));
  switch_elements_Calculator U_C
       (.\A0_reg[11]_0 (a0),
        .\B1_reg[11]_0 (b1),
        .D(a1),
        .FREQ(FREQ),
        .O(plusOp18),
        .Q(sh),
        .\a0d_reg[11] (st),
        .clk_i(clk_i),
        .\d1_4_reg[15] (z1i),
        .\d2_4_reg[15] (z2i),
        .\d3_4_reg[15] (z3i),
        .doii1(doii1),
        .out(out),
        .rst_i(rst_i),
        .\shii_reg[0]_0 (U_C_n_40),
        .\t3z3_reg[18] (p_1_in__0),
        .\z1d1_reg[15] (Q),
        .\z1d1_reg[15]_0 (tt1),
        .\z1d1_reg[15]_1 (d1_4),
        .\z1d1_reg[15]_2 (d78_1),
        .\z2d1_reg[15] (d56_2),
        .\z2d1_reg[15]_0 ({DZ2_78_n_0,DZ2_78_n_1,DZ2_78_n_2,DZ2_78_n_3,DZ2_78_n_4,DZ2_78_n_5,DZ2_78_n_6,DZ2_78_n_7,DZ2_78_n_8,DZ2_78_n_9,DZ2_78_n_10,DZ2_78_n_11,DZ2_78_n_12,DZ2_78_n_13,DZ2_78_n_14,DZ2_78_n_15}),
        .\z2d1_reg[15]_1 (d2_4),
        .\z2d1_reg[15]_2 (d78_2),
        .\z3d1_reg[15] (d56_3),
        .\z3d1_reg[15]_0 ({DZ3_78_n_1,DZ3_78_n_2,DZ3_78_n_3,DZ3_78_n_4,DZ3_78_n_5,DZ3_78_n_6,DZ3_78_n_7,DZ3_78_n_8,DZ3_78_n_9,DZ3_78_n_10,DZ3_78_n_11,DZ3_78_n_12,DZ3_78_n_13,DZ3_78_n_14,DZ3_78_n_15,DZ3_78_n_16}),
        .\z3d1_reg[15]_1 (d3_4),
        .\z3d1_reg[15]_2 (d78_3));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[0]),
        .Q(a0d[0]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[10]),
        .Q(a0d[10]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[11]),
        .Q(a0d[11]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[1]),
        .Q(a0d[1]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[2]),
        .Q(a0d[2]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[3]),
        .Q(a0d[3]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[4]),
        .Q(a0d[4]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[5]),
        .Q(a0d[5]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[6]),
        .Q(a0d[6]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[7]),
        .Q(a0d[7]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[8]),
        .Q(a0d[8]));
  FDCE #(
    .INIT(1'b0)) 
    \a0d_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a0[9]),
        .Q(a0d[9]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[0]),
        .Q(a1d[0]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[10]),
        .Q(a1d[10]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[11]),
        .Q(a1d[11]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[1]),
        .Q(a1d[1]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[2]),
        .Q(a1d[2]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[3]),
        .Q(a1d[3]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[4]),
        .Q(a1d[4]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[5]),
        .Q(a1d[5]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[6]),
        .Q(a1d[6]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[7]),
        .Q(a1d[7]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[8]),
        .Q(a1d[8]));
  FDCE #(
    .INIT(1'b0)) 
    \a1d_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(a1[9]),
        .Q(a1d[9]));
  LUT3 #(
    .INIT(8'h28)) 
    activity_blocks_c_9_i_1
       (.I0(st[2]),
        .I1(st[0]),
        .I2(st[1]),
        .O(d4_30));
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__72
       (.I0(\d4_40_reg[15]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__72_n_0));
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__73
       (.I0(\d4_40_reg[14]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__73_n_0));
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__74
       (.I0(\d4_40_reg[13]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__74_n_0));
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__75
       (.I0(\d4_40_reg[12]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__75_n_0));
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__76
       (.I0(\d4_40_reg[11]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__76_n_0));
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__77
       (.I0(\d4_40_reg[10]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__77_n_0));
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__78
       (.I0(\d4_40_reg[9]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__78_n_0));
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__79
       (.I0(\d4_40_reg[8]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__79_n_0));
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__80
       (.I0(\d4_40_reg[7]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__80_n_0));
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__81
       (.I0(\d4_40_reg[6]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__81_n_0));
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__82
       (.I0(\d4_40_reg[5]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__82_n_0));
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__83
       (.I0(\d4_40_reg[4]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__83_n_0));
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__84
       (.I0(\d4_40_reg[3]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__84_n_0));
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__85
       (.I0(\d4_40_reg[2]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__85_n_0));
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__86
       (.I0(\d4_40_reg[1]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__86_n_0));
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__87
       (.I0(\d4_40_reg[0]_activity_blocks_c_11_n_0 ),
        .I1(\d4_4_reg[15]_0 ),
        .O(activity_blocks_gate__87_n_0));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[0]),
        .Q(b1d[0]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[10]),
        .Q(b1d[10]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[11]),
        .Q(b1d[11]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[1]),
        .Q(b1d[1]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[2]),
        .Q(b1d[2]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[3]),
        .Q(b1d[3]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[4]),
        .Q(b1d[4]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[5]),
        .Q(b1d[5]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[6]),
        .Q(b1d[6]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[7]),
        .Q(b1d[7]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[8]),
        .Q(b1d[8]));
  FDCE #(
    .INIT(1'b0)) 
    \b1d_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(b1[9]),
        .Q(b1d[9]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[0] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[0]),
        .Q(d1_3[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[10] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[10]),
        .Q(d1_3[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[11] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[11]),
        .Q(d1_3[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[12] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[12]),
        .Q(d1_3[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[13] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[13]),
        .Q(d1_3[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[14] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[14]),
        .Q(d1_3[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[15] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[15]),
        .Q(d1_3[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[1] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[1]),
        .Q(d1_3[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[2] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[2]),
        .Q(d1_3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[3] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[3]),
        .Q(d1_3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[4] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[4]),
        .Q(d1_3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[5] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[5]),
        .Q(d1_3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[6] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[6]),
        .Q(d1_3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[7] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[7]),
        .Q(d1_3[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[8] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[8]),
        .Q(d1_3[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_3_reg[9] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(tt1[9]),
        .Q(d1_3[9]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[0] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[0]),
        .Q(d1_4[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[10] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[10]),
        .Q(d1_4[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[11] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[11]),
        .Q(d1_4[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[12] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[12]),
        .Q(d1_4[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[13] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[13]),
        .Q(d1_4[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[14] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[14]),
        .Q(d1_4[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[15] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[15]),
        .Q(d1_4[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[1] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[1]),
        .Q(d1_4[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[2] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[2]),
        .Q(d1_4[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[3] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[3]),
        .Q(d1_4[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[4] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[4]),
        .Q(d1_4[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[5] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[5]),
        .Q(d1_4[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[6] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[6]),
        .Q(d1_4[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[7] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[7]),
        .Q(d1_4[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[8] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[8]),
        .Q(d1_4[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d1_4_reg[9] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d1_3[9]),
        .Q(d1_4[9]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[0] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_15),
        .Q(d2_3[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[10] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_5),
        .Q(d2_3[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[11] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_4),
        .Q(d2_3[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[12] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_3),
        .Q(d2_3[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[13] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_2),
        .Q(d2_3[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[14] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_1),
        .Q(d2_3[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[15] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_0),
        .Q(d2_3[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[1] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_14),
        .Q(d2_3[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[2] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_13),
        .Q(d2_3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[3] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_12),
        .Q(d2_3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[4] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_11),
        .Q(d2_3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[5] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_10),
        .Q(d2_3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[6] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_9),
        .Q(d2_3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[7] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_8),
        .Q(d2_3[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[8] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_7),
        .Q(d2_3[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_3_reg[9] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ2_78_n_6),
        .Q(d2_3[9]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[0] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[0]),
        .Q(d2_4[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[10] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[10]),
        .Q(d2_4[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[11] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[11]),
        .Q(d2_4[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[12] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[12]),
        .Q(d2_4[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[13] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[13]),
        .Q(d2_4[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[14] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[14]),
        .Q(d2_4[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[15] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[15]),
        .Q(d2_4[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[1] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[1]),
        .Q(d2_4[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[2] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[2]),
        .Q(d2_4[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[3] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[3]),
        .Q(d2_4[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[4] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[4]),
        .Q(d2_4[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[5] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[5]),
        .Q(d2_4[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[6] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[6]),
        .Q(d2_4[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[7] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[7]),
        .Q(d2_4[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[8] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[8]),
        .Q(d2_4[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d2_4_reg[9] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d2_3[9]),
        .Q(d2_4[9]));
  LUT2 #(
    .INIT(4'h1)) 
    \d3_3[15]_i_1 
       (.I0(st[1]),
        .I1(st[2]),
        .O(a14));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[0] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_16),
        .Q(d3_3[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[10] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_6),
        .Q(d3_3[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[11] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_5),
        .Q(d3_3[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[12] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_4),
        .Q(d3_3[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[13] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_3),
        .Q(d3_3[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[14] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_2),
        .Q(d3_3[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[15] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_1),
        .Q(d3_3[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[1] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_15),
        .Q(d3_3[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[2] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_14),
        .Q(d3_3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[3] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_13),
        .Q(d3_3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[4] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_12),
        .Q(d3_3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[5] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_11),
        .Q(d3_3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[6] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_10),
        .Q(d3_3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[7] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_9),
        .Q(d3_3[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[8] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_8),
        .Q(d3_3[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_3_reg[9] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(DZ3_78_n_7),
        .Q(d3_3[9]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[0] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[0]),
        .Q(d3_4[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[10] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[10]),
        .Q(d3_4[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[11] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[11]),
        .Q(d3_4[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[12] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[12]),
        .Q(d3_4[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[13] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[13]),
        .Q(d3_4[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[14] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[14]),
        .Q(d3_4[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[15] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[15]),
        .Q(d3_4[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[1] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[1]),
        .Q(d3_4[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[2] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[2]),
        .Q(d3_4[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[3] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[3]),
        .Q(d3_4[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[4] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[4]),
        .Q(d3_4[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[5] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[5]),
        .Q(d3_4[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[6] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[6]),
        .Q(d3_4[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[7] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[7]),
        .Q(d3_4[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[8] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[8]),
        .Q(d3_4[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d3_4_reg[9] 
       (.C(clk_i),
        .CE(a14),
        .CLR(rst_i),
        .D(d3_3[9]),
        .Q(d3_4[9]));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[0]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[0]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[0]),
        .Q(\d4_3_reg[0]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[10]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[10]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[10]),
        .Q(\d4_3_reg[10]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[11]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[11]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[11]),
        .Q(\d4_3_reg[11]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[12]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[12]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[12]),
        .Q(\d4_3_reg[12]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[13]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[13]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[13]),
        .Q(\d4_3_reg[13]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[14]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[14]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[14]),
        .Q(\d4_3_reg[14]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[15]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[15]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[15]),
        .Q(\d4_3_reg[15]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[1]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[1]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[1]),
        .Q(\d4_3_reg[1]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[2]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[2]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[2]),
        .Q(\d4_3_reg[2]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[3]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[3]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[3]),
        .Q(\d4_3_reg[3]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[4]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[4]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[4]),
        .Q(\d4_3_reg[4]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[5]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[5]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[5]),
        .Q(\d4_3_reg[5]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[6]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[6]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[6]),
        .Q(\d4_3_reg[6]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[7]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[7]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[7]),
        .Q(\d4_3_reg[7]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[8]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[8]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[8]),
        .Q(\d4_3_reg[8]_srl2_activity_blocks_c_10_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutG/d4_3_reg " *) 
  (* srl_name = "\activity_blocks[0].dutG/d4_3_reg[9]_srl2_activity_blocks_c_10 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \d4_3_reg[9]_srl2_activity_blocks_c_10 
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(d4_30),
        .CLK(clk_i),
        .D(dd2[9]),
        .Q(\d4_3_reg[9]_srl2_activity_blocks_c_10_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[0]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[0]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[0]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[10]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[10]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[10]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[11]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[11]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[11]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[12]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[12]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[12]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[13]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[13]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[13]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[14]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[14]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[14]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[15]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[15]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[15]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[1]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[1]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[1]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[2]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[2]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[2]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[3]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[3]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[3]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[4]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[4]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[4]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[5]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[5]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[5]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[6]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[6]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[6]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[7]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[7]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[7]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[8]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[8]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[8]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \d4_40_reg[9]_activity_blocks_c_11 
       (.C(clk_i),
        .CE(d4_30),
        .D(\d4_3_reg[9]_srl2_activity_blocks_c_10_n_0 ),
        .Q(\d4_40_reg[9]_activity_blocks_c_11_n_0 ),
        .R(1'b0));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[0] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__87_n_0),
        .Q(d4_4[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[10] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__77_n_0),
        .Q(d4_4[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[11] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__76_n_0),
        .Q(d4_4[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[12] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__75_n_0),
        .Q(d4_4[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[13] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__74_n_0),
        .Q(d4_4[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[14] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__73_n_0),
        .Q(d4_4[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[15] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__72_n_0),
        .Q(d4_4[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[1] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__86_n_0),
        .Q(d4_4[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[2] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__85_n_0),
        .Q(d4_4[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[3] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__84_n_0),
        .Q(d4_4[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[4] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__83_n_0),
        .Q(d4_4[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[5] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__82_n_0),
        .Q(d4_4[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[6] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__81_n_0),
        .Q(d4_4[6]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[7] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__80_n_0),
        .Q(d4_4[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[8] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__79_n_0),
        .Q(d4_4[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d4_4_reg[9] 
       (.C(clk_i),
        .CE(d4_30),
        .CLR(rst_i),
        .D(activity_blocks_gate__78_n_0),
        .Q(d4_4[9]));
  LUT4 #(
    .INIT(16'h0008)) 
    \d_z2[20]_i_2 
       (.I0(did[15]),
        .I1(st[0]),
        .I2(st[1]),
        .I3(st[2]),
        .O(\d_z2[20]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \d_z2[20]_i_3 
       (.I0(did[14]),
        .I1(st[0]),
        .I2(st[1]),
        .I3(st[2]),
        .O(\d_z2[20]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \d_z2[20]_i_4 
       (.I0(st[2]),
        .I1(st[1]),
        .I2(st[0]),
        .I3(did[15]),
        .O(\d_z2[20]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \d_z2[20]_i_5 
       (.I0(st[2]),
        .I1(st[1]),
        .I2(st[0]),
        .I3(did[15]),
        .O(\d_z2[20]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \d_z2[20]_i_6 
       (.I0(st[2]),
        .I1(st[1]),
        .I2(st[0]),
        .I3(did[14]),
        .O(\d_z2[20]_i_6_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[10]),
        .Q(A[7]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[11]),
        .Q(A[8]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[12]),
        .Q(A[9]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[13]),
        .Q(A[10]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[14]),
        .Q(A[11]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[15]),
        .Q(A[12]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[16]),
        .Q(A[13]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[17]),
        .Q(A[14]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[18]),
        .Q(A[15]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[20]),
        .Q(A[17]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[3]),
        .Q(A[0]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[4]),
        .Q(A[1]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[5]),
        .Q(A[2]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[6]),
        .Q(A[3]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[7]),
        .Q(A[4]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[8]),
        .Q(A[5]));
  FDCE #(
    .INIT(1'b0)) 
    \d_z2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(minusOp[9]),
        .Q(A[6]));
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \dd1[16]_i_1 
       (.I0(did[14]),
        .I1(st[0]),
        .I2(st[1]),
        .I3(st[2]),
        .O(dii[16]));
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \dd1[18]_i_1 
       (.I0(did[15]),
        .I1(st[0]),
        .I2(st[1]),
        .I3(st[2]),
        .O(dii[18]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[0]),
        .Q(dd1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[10]),
        .Q(dd1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[11]),
        .Q(dd1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[12]),
        .Q(dd1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[13]),
        .Q(dd1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[14]),
        .Q(dd1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[15]),
        .Q(dd1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[16]),
        .Q(dd1[16]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[18]),
        .Q(dd1[18]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[1]),
        .Q(dd1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[2]),
        .Q(dd1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[3]),
        .Q(dd1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[4]),
        .Q(dd1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[5]),
        .Q(dd1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[6]),
        .Q(dd1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[7]),
        .Q(dd1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[8]),
        .Q(dd1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \dd1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dii[9]),
        .Q(dd1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[0]),
        .Q(dd2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[10]),
        .Q(dd2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[11]),
        .Q(dd2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[12]),
        .Q(dd2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[13]),
        .Q(dd2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[14]),
        .Q(dd2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[15]),
        .Q(dd2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[16]),
        .Q(dd2__0[16]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[18]),
        .Q(dd2__0[18]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[1]),
        .Q(dd2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[2]),
        .Q(dd2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[3]),
        .Q(dd2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[4]),
        .Q(dd2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[5]),
        .Q(dd2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[6]),
        .Q(dd2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[7]),
        .Q(dd2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[8]),
        .Q(dd2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \dd2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(dd1[9]),
        .Q(dd2[9]));
  LUT3 #(
    .INIT(8'h01)) 
    \did[15]_i_1 
       (.I0(st[1]),
        .I1(st[2]),
        .I2(st[0]),
        .O(\did[15]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[0] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[0]),
        .Q(did[0]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[10] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[10]),
        .Q(did[10]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[11] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[11]),
        .Q(did[11]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[12] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[12]),
        .Q(did[12]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[13] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[13]),
        .Q(did[13]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[14] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[14]),
        .Q(did[14]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[15] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[15]),
        .Q(did[15]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[1] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[1]),
        .Q(did[1]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[2] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[2]),
        .Q(did[2]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[3] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[3]),
        .Q(did[3]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[4] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[4]),
        .Q(did[4]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[5] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[5]),
        .Q(did[5]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[6] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[6]),
        .Q(did[6]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[7] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[7]),
        .Q(did[7]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[8] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[8]),
        .Q(did[8]));
  FDCE #(
    .INIT(1'b0)) 
    \did_reg[9] 
       (.C(clk_i),
        .CE(\did[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(DI[9]),
        .Q(did[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \st[0]_i_1__0 
       (.I0(st[0]),
        .O(\st[0]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \st[1]_i_1__0 
       (.I0(st[0]),
        .I1(st[1]),
        .O(\st[1]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \st[2]_i_1__0 
       (.I0(st[1]),
        .I1(st[0]),
        .I2(st[2]),
        .O(\st[2]_i_1__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\st[0]_i_1__0_n_0 ),
        .Q(st[0]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\st[1]_i_1__0_n_0 ),
        .Q(st[1]));
  FDCE #(
    .INIT(1'b0)) 
    \st_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\st[2]_i_1__0_n_0 ),
        .Q(st[2]));
  (* ACASCREG = "0" *) 
  (* ADREG = "1" *) 
  (* ALUMODEREG = "0" *) 
  (* AMULTSEL = "A" *) 
  (* AREG = "0" *) 
  (* AUTORESET_PATDET = "NO_RESET" *) 
  (* AUTORESET_PRIORITY = "RESET" *) 
  (* A_INPUT = "DIRECT" *) 
  (* BCASCREG = "0" *) 
  (* BMULTSEL = "B" *) 
  (* BREG = "0" *) 
  (* B_INPUT = "DIRECT" *) 
  (* CARRYINREG = "0" *) 
  (* CARRYINSELREG = "0" *) 
  (* CREG = "0" *) 
  (* DREG = "1" *) 
  (* INMODEREG = "0" *) 
  (* MASK = "48'h3FFFFFFFFFFF" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  (* MREG = "0" *) 
  (* OPMODEREG = "0" *) 
  (* PATTERN = "48'h000000000000" *) 
  (* PREADDINSEL = "A" *) 
  (* PREG = "1" *) 
  (* RND = "48'h000000000000" *) 
  (* SEL_MASK = "MASK" *) 
  (* SEL_PATTERN = "PATTERN" *) 
  (* USE_MULT = "MULTIPLY" *) 
  (* USE_PATTERN_DETECT = "NO_PATDET" *) 
  (* USE_SIMD = "ONE48" *) 
  (* USE_WIDEXOR = "FALSE" *) 
  (* XORSIMD = "XOR24_48_96" *) 
  DSP48E2_UNIQ_BASE_ t1_reg
       (.A({tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1[21],tt2_z1}),
        .ACIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .ACOUT(NLW_t1_reg_ACOUT_UNCONNECTED[29:0]),
        .ALUMODE({1'b0,1'b0,1'b0,1'b0}),
        .B({a1d[11],a1d[11],a1d[11],a1d[11],a1d[11],a1d[11],a1d}),
        .BCIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .BCOUT(NLW_t1_reg_BCOUT_UNCONNECTED[17:0]),
        .C({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CARRYCASCIN(1'b0),
        .CARRYCASCOUT(NLW_t1_reg_CARRYCASCOUT_UNCONNECTED),
        .CARRYIN(1'b0),
        .CARRYINSEL({1'b0,1'b0,1'b0}),
        .CARRYOUT(NLW_t1_reg_CARRYOUT_UNCONNECTED[3:0]),
        .CEA1(1'b0),
        .CEA2(1'b0),
        .CEAD(1'b0),
        .CEALUMODE(1'b0),
        .CEB1(1'b0),
        .CEB2(1'b0),
        .CEC(1'b0),
        .CECARRYIN(1'b0),
        .CECTRL(1'b0),
        .CED(1'b0),
        .CEINMODE(1'b0),
        .CEM(1'b0),
        .CEP(1'b1),
        .CLK(clk_i),
        .D({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .INMODE({1'b0,1'b0,1'b0,1'b0,1'b0}),
        .MULTSIGNIN(1'b0),
        .MULTSIGNOUT(NLW_t1_reg_MULTSIGNOUT_UNCONNECTED),
        .OPMODE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}),
        .OVERFLOW(NLW_t1_reg_OVERFLOW_UNCONNECTED),
        .P({NLW_t1_reg_P_UNCONNECTED[47:29],t1_reg_n_77,t1_reg_n_78,t1_reg_n_79,t1_reg_n_80,t1_reg_n_81,t1_reg_n_82,t1_reg_n_83,t1_reg_n_84,t1_reg_n_85,t1_reg_n_86,t1_reg_n_87,t1_reg_n_88,t1_reg_n_89,t1_reg_n_90,t1_reg_n_91,t1_reg_n_92,t1_reg_n_93,t1_reg_n_94,t1_reg_n_95,t1_reg_n_96,t1_reg_n_97,t1_reg_n_98,t1_reg_n_99,t1_reg_n_100,t1_reg_n_101,t1_reg_n_102,t1_reg_n_103,t1_reg_n_104,t1_reg_n_105}),
        .PATTERNBDETECT(NLW_t1_reg_PATTERNBDETECT_UNCONNECTED),
        .PATTERNDETECT(NLW_t1_reg_PATTERNDETECT_UNCONNECTED),
        .PCIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .PCOUT(NLW_t1_reg_PCOUT_UNCONNECTED[47:0]),
        .RSTA(1'b0),
        .RSTALLCARRYIN(1'b0),
        .RSTALUMODE(1'b0),
        .RSTB(1'b0),
        .RSTC(1'b0),
        .RSTCTRL(1'b0),
        .RSTD(1'b0),
        .RSTINMODE(1'b0),
        .RSTM(1'b0),
        .RSTP(1'b0),
        .UNDERFLOW(NLW_t1_reg_UNDERFLOW_UNCONNECTED),
        .XOROUT(NLW_t1_reg_XOROUT_UNCONNECTED[7:0]));
  (* ACASCREG = "0" *) 
  (* ADREG = "1" *) 
  (* ALUMODEREG = "0" *) 
  (* AMULTSEL = "A" *) 
  (* AREG = "0" *) 
  (* AUTORESET_PATDET = "NO_RESET" *) 
  (* AUTORESET_PRIORITY = "RESET" *) 
  (* A_INPUT = "DIRECT" *) 
  (* BCASCREG = "0" *) 
  (* BMULTSEL = "B" *) 
  (* BREG = "0" *) 
  (* B_INPUT = "DIRECT" *) 
  (* CARRYINREG = "0" *) 
  (* CARRYINSELREG = "0" *) 
  (* CREG = "0" *) 
  (* DREG = "1" *) 
  (* INMODEREG = "0" *) 
  (* MASK = "48'h3FFFFFFFFFFF" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  (* MREG = "0" *) 
  (* OPMODEREG = "0" *) 
  (* PATTERN = "48'h000000000000" *) 
  (* PREADDINSEL = "A" *) 
  (* PREG = "1" *) 
  (* RND = "48'h000000000000" *) 
  (* SEL_MASK = "MASK" *) 
  (* SEL_PATTERN = "PATTERN" *) 
  (* USE_MULT = "MULTIPLY" *) 
  (* USE_PATTERN_DETECT = "NO_PATDET" *) 
  (* USE_SIMD = "ONE48" *) 
  (* USE_WIDEXOR = "FALSE" *) 
  (* XORSIMD = "XOR24_48_96" *) 
  DSP48E2_HD32740 t2_reg
       (.A({A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[17],A[15:0]}),
        .ACIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .ACOUT(NLW_t2_reg_ACOUT_UNCONNECTED[29:0]),
        .ALUMODE({1'b0,1'b0,1'b0,1'b0}),
        .B({b1d[11],b1d[11],b1d[11],b1d[11],b1d[11],b1d[11],b1d}),
        .BCIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .BCOUT(NLW_t2_reg_BCOUT_UNCONNECTED[17:0]),
        .C({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CARRYCASCIN(1'b0),
        .CARRYCASCOUT(NLW_t2_reg_CARRYCASCOUT_UNCONNECTED),
        .CARRYIN(1'b0),
        .CARRYINSEL({1'b0,1'b0,1'b0}),
        .CARRYOUT(NLW_t2_reg_CARRYOUT_UNCONNECTED[3:0]),
        .CEA1(1'b0),
        .CEA2(1'b0),
        .CEAD(1'b0),
        .CEALUMODE(1'b0),
        .CEB1(1'b0),
        .CEB2(1'b0),
        .CEC(1'b0),
        .CECARRYIN(1'b0),
        .CECTRL(1'b0),
        .CED(1'b0),
        .CEINMODE(1'b0),
        .CEM(1'b0),
        .CEP(1'b1),
        .CLK(clk_i),
        .D({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .INMODE({1'b0,1'b0,1'b0,1'b0,1'b0}),
        .MULTSIGNIN(1'b0),
        .MULTSIGNOUT(NLW_t2_reg_MULTSIGNOUT_UNCONNECTED),
        .OPMODE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}),
        .OVERFLOW(NLW_t2_reg_OVERFLOW_UNCONNECTED),
        .P({NLW_t2_reg_P_UNCONNECTED[47:29],t2_reg_n_77,R,t2_reg_n_98,t2_reg_n_99,t2_reg_n_100,t2_reg_n_101,t2_reg_n_102,t2_reg_n_103,t2_reg_n_104,t2_reg_n_105}),
        .PATTERNBDETECT(NLW_t2_reg_PATTERNBDETECT_UNCONNECTED),
        .PATTERNDETECT(NLW_t2_reg_PATTERNDETECT_UNCONNECTED),
        .PCIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .PCOUT(NLW_t2_reg_PCOUT_UNCONNECTED[47:0]),
        .RSTA(1'b0),
        .RSTALLCARRYIN(1'b0),
        .RSTALUMODE(1'b0),
        .RSTB(1'b0),
        .RSTC(1'b0),
        .RSTCTRL(1'b0),
        .RSTD(1'b0),
        .RSTINMODE(1'b0),
        .RSTM(1'b0),
        .RSTP(1'b0),
        .UNDERFLOW(NLW_t2_reg_UNDERFLOW_UNCONNECTED),
        .XOROUT(NLW_t2_reg_XOROUT_UNCONNECTED[7:0]));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_2 
       (.I0(z2d2[15]),
        .I1(R[15]),
        .O(\t2z2[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_3 
       (.I0(z2d2[14]),
        .I1(R[14]),
        .O(\t2z2[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_4 
       (.I0(z2d2[13]),
        .I1(R[13]),
        .O(\t2z2[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_5 
       (.I0(z2d2[12]),
        .I1(R[12]),
        .O(\t2z2[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_6 
       (.I0(z2d2[11]),
        .I1(R[11]),
        .O(\t2z2[15]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_7 
       (.I0(z2d2[10]),
        .I1(R[10]),
        .O(\t2z2[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_8 
       (.I0(z2d2[9]),
        .I1(R[9]),
        .O(\t2z2[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[15]_i_9 
       (.I0(z2d2[8]),
        .I1(R[8]),
        .O(\t2z2[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_2 
       (.I0(z2d2[7]),
        .I1(R[7]),
        .O(\t2z2[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_3 
       (.I0(z2d2[6]),
        .I1(R[6]),
        .O(\t2z2[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_4 
       (.I0(z2d2[5]),
        .I1(R[5]),
        .O(\t2z2[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_5 
       (.I0(z2d2[4]),
        .I1(R[4]),
        .O(\t2z2[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_6 
       (.I0(z2d2[3]),
        .I1(R[3]),
        .O(\t2z2[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_7 
       (.I0(z2d2[2]),
        .I1(R[2]),
        .O(\t2z2[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_8 
       (.I0(z2d2[1]),
        .I1(R[1]),
        .O(\t2z2[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t2z2[7]_i_9 
       (.I0(z2d2[0]),
        .I1(R[0]),
        .O(\t2z2[7]_i_9_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[0]),
        .Q(t2z2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[10]),
        .Q(t2z2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[11]),
        .Q(t2z2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[12]),
        .Q(t2z2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[13]),
        .Q(t2z2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[14]),
        .Q(t2z2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[15]),
        .Q(t2z2[15]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t2z2_reg[15]_i_1 
       (.CI(\t2z2_reg[7]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\t2z2_reg[15]_i_1_n_0 ,\t2z2_reg[15]_i_1_n_1 ,\t2z2_reg[15]_i_1_n_2 ,\t2z2_reg[15]_i_1_n_3 ,\t2z2_reg[15]_i_1_n_4 ,\t2z2_reg[15]_i_1_n_5 ,\t2z2_reg[15]_i_1_n_6 ,\t2z2_reg[15]_i_1_n_7 }),
        .DI(z2d2[15:8]),
        .O(t2z2i[15:8]),
        .S({\t2z2[15]_i_2_n_0 ,\t2z2[15]_i_3_n_0 ,\t2z2[15]_i_4_n_0 ,\t2z2[15]_i_5_n_0 ,\t2z2[15]_i_6_n_0 ,\t2z2[15]_i_7_n_0 ,\t2z2[15]_i_8_n_0 ,\t2z2[15]_i_9_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[16]),
        .Q(t2z2[16]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[17]),
        .Q(t2z2[17]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[18]),
        .Q(t2z2[18]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[19]),
        .Q(t2z2[19]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t2z2_reg[19]_i_1 
       (.CI(\t2z2_reg[15]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_t2z2_reg[19]_i_1_CO_UNCONNECTED [7:3],\t2z2_reg[19]_i_1_n_5 ,\t2z2_reg[19]_i_1_n_6 ,\t2z2_reg[19]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_t2z2_reg[19]_i_1_O_UNCONNECTED [7:4],t2z2i[19:16]}),
        .S({1'b0,1'b0,1'b0,1'b0,R[19:16]}));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[1]),
        .Q(t2z2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[2]),
        .Q(t2z2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[3]),
        .Q(t2z2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[4]),
        .Q(t2z2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[5]),
        .Q(t2z2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[6]),
        .Q(t2z2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[7]),
        .Q(t2z2[7]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t2z2_reg[7]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\t2z2_reg[7]_i_1_n_0 ,\t2z2_reg[7]_i_1_n_1 ,\t2z2_reg[7]_i_1_n_2 ,\t2z2_reg[7]_i_1_n_3 ,\t2z2_reg[7]_i_1_n_4 ,\t2z2_reg[7]_i_1_n_5 ,\t2z2_reg[7]_i_1_n_6 ,\t2z2_reg[7]_i_1_n_7 }),
        .DI(z2d2[7:0]),
        .O(t2z2i[7:0]),
        .S({\t2z2[7]_i_2_n_0 ,\t2z2[7]_i_3_n_0 ,\t2z2[7]_i_4_n_0 ,\t2z2[7]_i_5_n_0 ,\t2z2[7]_i_6_n_0 ,\t2z2[7]_i_7_n_0 ,\t2z2[7]_i_8_n_0 ,\t2z2[7]_i_9_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[8]),
        .Q(t2z2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2i[9]),
        .Q(t2z2[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \t2z2_z3[19]_i_2 
       (.I0(t2z2[19]),
        .O(\t2z2_z3[19]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \t2z2_z3[19]_i_3 
       (.I0(t2z2[18]),
        .O(\t2z2_z3[19]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \t2z2_z3[19]_i_4 
       (.I0(t2z2[17]),
        .O(\t2z2_z3[19]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \t2z2_z3[19]_i_5 
       (.I0(t2z2[16]),
        .O(\t2z2_z3[19]_i_5_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_25),
        .Q(t2z2_z3[10]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_24),
        .Q(t2z2_z3[11]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_23),
        .Q(t2z2_z3[12]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_22),
        .Q(t2z2_z3[13]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_21),
        .Q(t2z2_z3[14]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_20),
        .Q(t2z2_z3[15]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_19),
        .Q(t2z2_z3[16]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_18),
        .Q(t2z2_z3[17]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_17),
        .Q(t2z2_z3[18]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_16),
        .Q(t2z2_z3[19]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_33),
        .Q(t2z2_z3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_32),
        .Q(t2z2_z3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_31),
        .Q(t2z2_z3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_30),
        .Q(t2z2_z3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_29),
        .Q(t2z2_z3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_28),
        .Q(t2z2_z3[7]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_27),
        .Q(t2z2_z3[8]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2_z3_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ3_n_26),
        .Q(t2z2_z3[9]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[0]),
        .Q(t2z2d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[10]),
        .Q(t2z2d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[11]),
        .Q(t2z2d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[12]),
        .Q(t2z2d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[13]),
        .Q(t2z2d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[14]),
        .Q(t2z2d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[15]),
        .Q(t2z2d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[1]),
        .Q(t2z2d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[2]),
        .Q(t2z2d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[3]),
        .Q(t2z2d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[4]),
        .Q(t2z2d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[5]),
        .Q(t2z2d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[6]),
        .Q(t2z2d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[7]),
        .Q(t2z2d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[8]),
        .Q(t2z2d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2[9]),
        .Q(t2z2d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[0]),
        .Q(t2z2d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[10]),
        .Q(t2z2d2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[11]),
        .Q(t2z2d2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[12]),
        .Q(t2z2d2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[13]),
        .Q(t2z2d2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[14]),
        .Q(t2z2d2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[15]),
        .Q(t2z2d2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[1]),
        .Q(t2z2d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[2]),
        .Q(t2z2d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[3]),
        .Q(t2z2d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[4]),
        .Q(t2z2d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[5]),
        .Q(t2z2d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[6]),
        .Q(t2z2d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[7]),
        .Q(t2z2d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[8]),
        .Q(t2z2d2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \t2z2d2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(t2z2d1[9]),
        .Q(t2z2d2[9]));
  (* ACASCREG = "0" *) 
  (* ADREG = "1" *) 
  (* ALUMODEREG = "0" *) 
  (* AMULTSEL = "A" *) 
  (* AREG = "0" *) 
  (* AUTORESET_PATDET = "NO_RESET" *) 
  (* AUTORESET_PRIORITY = "RESET" *) 
  (* A_INPUT = "DIRECT" *) 
  (* BCASCREG = "0" *) 
  (* BMULTSEL = "B" *) 
  (* BREG = "0" *) 
  (* B_INPUT = "DIRECT" *) 
  (* CARRYINREG = "0" *) 
  (* CARRYINSELREG = "0" *) 
  (* CREG = "0" *) 
  (* DREG = "1" *) 
  (* INMODEREG = "0" *) 
  (* MASK = "48'h3FFFFFFFFFFF" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  (* MREG = "0" *) 
  (* OPMODEREG = "0" *) 
  (* PATTERN = "48'h000000000000" *) 
  (* PREADDINSEL = "A" *) 
  (* PREG = "1" *) 
  (* RND = "48'h000000000000" *) 
  (* SEL_MASK = "MASK" *) 
  (* SEL_PATTERN = "PATTERN" *) 
  (* USE_MULT = "MULTIPLY" *) 
  (* USE_PATTERN_DETECT = "NO_PATDET" *) 
  (* USE_SIMD = "ONE48" *) 
  (* USE_WIDEXOR = "FALSE" *) 
  (* XORSIMD = "XOR24_48_96" *) 
  DSP48E2_HD32741 t3_reg
       (.A({t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3[19],t2z2_z3}),
        .ACIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .ACOUT(NLW_t3_reg_ACOUT_UNCONNECTED[29:0]),
        .ALUMODE({1'b0,1'b0,1'b0,1'b0}),
        .B({a0d[11],a0d[11],a0d[11],a0d[11],a0d[11],a0d[11],a0d}),
        .BCIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .BCOUT(NLW_t3_reg_BCOUT_UNCONNECTED[17:0]),
        .C({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CARRYCASCIN(1'b0),
        .CARRYCASCOUT(NLW_t3_reg_CARRYCASCOUT_UNCONNECTED),
        .CARRYIN(1'b0),
        .CARRYINSEL({1'b0,1'b0,1'b0}),
        .CARRYOUT(NLW_t3_reg_CARRYOUT_UNCONNECTED[3:0]),
        .CEA1(1'b0),
        .CEA2(1'b0),
        .CEAD(1'b0),
        .CEALUMODE(1'b0),
        .CEB1(1'b0),
        .CEB2(1'b0),
        .CEC(1'b0),
        .CECARRYIN(1'b0),
        .CECTRL(1'b0),
        .CED(1'b0),
        .CEINMODE(1'b0),
        .CEM(1'b0),
        .CEP(1'b1),
        .CLK(clk_i),
        .D({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .INMODE({1'b0,1'b0,1'b0,1'b0,1'b0}),
        .MULTSIGNIN(1'b0),
        .MULTSIGNOUT(NLW_t3_reg_MULTSIGNOUT_UNCONNECTED),
        .OPMODE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}),
        .OVERFLOW(NLW_t3_reg_OVERFLOW_UNCONNECTED),
        .P({NLW_t3_reg_P_UNCONNECTED[47:29],t3_reg_n_77,L,t3_reg_n_97,t3_reg_n_98,t3_reg_n_99,t3_reg_n_100,t3_reg_n_101,t3_reg_n_102,t3_reg_n_103,t3_reg_n_104,t3_reg_n_105}),
        .PATTERNBDETECT(NLW_t3_reg_PATTERNBDETECT_UNCONNECTED),
        .PATTERNDETECT(NLW_t3_reg_PATTERNDETECT_UNCONNECTED),
        .PCIN({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .PCOUT(NLW_t3_reg_PCOUT_UNCONNECTED[47:0]),
        .RSTA(1'b0),
        .RSTALLCARRYIN(1'b0),
        .RSTALUMODE(1'b0),
        .RSTB(1'b0),
        .RSTC(1'b0),
        .RSTCTRL(1'b0),
        .RSTD(1'b0),
        .RSTINMODE(1'b0),
        .RSTM(1'b0),
        .RSTP(1'b0),
        .UNDERFLOW(NLW_t3_reg_UNDERFLOW_UNCONNECTED),
        .XOROUT(NLW_t3_reg_XOROUT_UNCONNECTED[7:0]));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_2 
       (.I0(z3d2[15]),
        .I1(L[24]),
        .O(\t3z3[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_3 
       (.I0(z3d2[14]),
        .I1(L[23]),
        .O(\t3z3[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_4 
       (.I0(z3d2[13]),
        .I1(L[22]),
        .O(\t3z3[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_5 
       (.I0(z3d2[12]),
        .I1(L[21]),
        .O(\t3z3[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_6 
       (.I0(z3d2[11]),
        .I1(L[20]),
        .O(\t3z3[15]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_7 
       (.I0(z3d2[10]),
        .I1(L[19]),
        .O(\t3z3[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_8 
       (.I0(z3d2[9]),
        .I1(L[18]),
        .O(\t3z3[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[15]_i_9 
       (.I0(z3d2[8]),
        .I1(L[17]),
        .O(\t3z3[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_2 
       (.I0(z3d2[7]),
        .I1(L[16]),
        .O(\t3z3[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_3 
       (.I0(z3d2[6]),
        .I1(L[15]),
        .O(\t3z3[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_4 
       (.I0(z3d2[5]),
        .I1(L[14]),
        .O(\t3z3[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_5 
       (.I0(z3d2[4]),
        .I1(L[13]),
        .O(\t3z3[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_6 
       (.I0(z3d2[3]),
        .I1(L[12]),
        .O(\t3z3[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_7 
       (.I0(z3d2[2]),
        .I1(L[11]),
        .O(\t3z3[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_8 
       (.I0(z3d2[1]),
        .I1(L[10]),
        .O(\t3z3[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \t3z3[7]_i_9 
       (.I0(z3d2[0]),
        .I1(L[9]),
        .O(\t3z3[7]_i_9_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[0]),
        .Q(t3z3[0]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[10]),
        .Q(t3z3[10]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[11]),
        .Q(t3z3[11]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[12]),
        .Q(t3z3[12]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[13]),
        .Q(t3z3[13]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[14]),
        .Q(t3z3[14]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[15]),
        .Q(t3z3[15]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t3z3_reg[15]_i_1 
       (.CI(\t3z3_reg[7]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\t3z3_reg[15]_i_1_n_0 ,\t3z3_reg[15]_i_1_n_1 ,\t3z3_reg[15]_i_1_n_2 ,\t3z3_reg[15]_i_1_n_3 ,\t3z3_reg[15]_i_1_n_4 ,\t3z3_reg[15]_i_1_n_5 ,\t3z3_reg[15]_i_1_n_6 ,\t3z3_reg[15]_i_1_n_7 }),
        .DI(z3d2[15:8]),
        .O(plusOp[15:8]),
        .S({\t3z3[15]_i_2_n_0 ,\t3z3[15]_i_3_n_0 ,\t3z3[15]_i_4_n_0 ,\t3z3[15]_i_5_n_0 ,\t3z3[15]_i_6_n_0 ,\t3z3[15]_i_7_n_0 ,\t3z3[15]_i_8_n_0 ,\t3z3[15]_i_9_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[16]),
        .Q(t3z3[16]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[17]),
        .Q(t3z3[17]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[18]),
        .Q(t3z3[18]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t3z3_reg[18]_i_1 
       (.CI(\t3z3_reg[15]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_t3z3_reg[18]_i_1_CO_UNCONNECTED [7:2],\t3z3_reg[18]_i_1_n_6 ,\t3z3_reg[18]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_t3z3_reg[18]_i_1_O_UNCONNECTED [7:3],plusOp[18:16]}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,L[27:25]}));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[1]),
        .Q(t3z3[1]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[2]),
        .Q(t3z3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[3]),
        .Q(t3z3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[4]),
        .Q(t3z3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[5]),
        .Q(t3z3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[6]),
        .Q(t3z3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[7]),
        .Q(t3z3[7]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \t3z3_reg[7]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\t3z3_reg[7]_i_1_n_0 ,\t3z3_reg[7]_i_1_n_1 ,\t3z3_reg[7]_i_1_n_2 ,\t3z3_reg[7]_i_1_n_3 ,\t3z3_reg[7]_i_1_n_4 ,\t3z3_reg[7]_i_1_n_5 ,\t3z3_reg[7]_i_1_n_6 ,\t3z3_reg[7]_i_1_n_7 }),
        .DI(z3d2[7:0]),
        .O(plusOp[7:0]),
        .S({\t3z3[7]_i_2_n_0 ,\t3z3[7]_i_3_n_0 ,\t3z3[7]_i_4_n_0 ,\t3z3[7]_i_5_n_0 ,\t3z3[7]_i_6_n_0 ,\t3z3[7]_i_7_n_0 ,\t3z3[7]_i_8_n_0 ,\t3z3[7]_i_9_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[8]),
        .Q(t3z3[8]));
  FDCE #(
    .INIT(1'b0)) 
    \t3z3_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(plusOp[9]),
        .Q(t3z3[9]));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_2 
       (.I0(dd2[15]),
        .I1(R[15]),
        .O(\tt2[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_3 
       (.I0(dd2[14]),
        .I1(R[14]),
        .O(\tt2[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_4 
       (.I0(dd2[13]),
        .I1(R[13]),
        .O(\tt2[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_5 
       (.I0(dd2[12]),
        .I1(R[12]),
        .O(\tt2[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_6 
       (.I0(dd2[11]),
        .I1(R[11]),
        .O(\tt2[15]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_7 
       (.I0(dd2[10]),
        .I1(R[10]),
        .O(\tt2[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_8 
       (.I0(dd2[9]),
        .I1(R[9]),
        .O(\tt2[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[15]_i_9 
       (.I0(dd2[8]),
        .I1(R[8]),
        .O(\tt2[15]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \tt2[20]_i_2 
       (.I0(R[18]),
        .O(\tt2[20]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2[20]_i_3 
       (.I0(R[19]),
        .I1(t2_reg_n_77),
        .O(\tt2[20]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \tt2[20]_i_4 
       (.I0(R[18]),
        .I1(R[19]),
        .O(\tt2[20]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[20]_i_5 
       (.I0(R[18]),
        .I1(dd2__0[18]),
        .O(\tt2[20]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[20]_i_6 
       (.I0(dd2__0[18]),
        .I1(R[17]),
        .O(\tt2[20]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[20]_i_7 
       (.I0(dd2__0[16]),
        .I1(R[16]),
        .O(\tt2[20]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_2 
       (.I0(dd2[7]),
        .I1(R[7]),
        .O(\tt2[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_3 
       (.I0(dd2[6]),
        .I1(R[6]),
        .O(\tt2[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_4 
       (.I0(dd2[5]),
        .I1(R[5]),
        .O(\tt2[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_5 
       (.I0(dd2[4]),
        .I1(R[4]),
        .O(\tt2[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_6 
       (.I0(dd2[3]),
        .I1(R[3]),
        .O(\tt2[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_7 
       (.I0(dd2[2]),
        .I1(R[2]),
        .O(\tt2[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_8 
       (.I0(dd2[1]),
        .I1(R[1]),
        .O(\tt2[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \tt2[7]_i_9 
       (.I0(dd2[0]),
        .I1(R[0]),
        .O(\tt2[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[0] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_15 ),
        .Q(tt2[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[10] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_13 ),
        .Q(tt2[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[11] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_12 ),
        .Q(tt2[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[12] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_11 ),
        .Q(tt2[12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[13] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_10 ),
        .Q(tt2[13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[14] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_9 ),
        .Q(tt2[14]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[15] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_8 ),
        .Q(tt2[15]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tt2_reg[15]_i_1 
       (.CI(\tt2_reg[7]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tt2_reg[15]_i_1_n_0 ,\tt2_reg[15]_i_1_n_1 ,\tt2_reg[15]_i_1_n_2 ,\tt2_reg[15]_i_1_n_3 ,\tt2_reg[15]_i_1_n_4 ,\tt2_reg[15]_i_1_n_5 ,\tt2_reg[15]_i_1_n_6 ,\tt2_reg[15]_i_1_n_7 }),
        .DI(dd2[15:8]),
        .O({\tt2_reg[15]_i_1_n_8 ,\tt2_reg[15]_i_1_n_9 ,\tt2_reg[15]_i_1_n_10 ,\tt2_reg[15]_i_1_n_11 ,\tt2_reg[15]_i_1_n_12 ,\tt2_reg[15]_i_1_n_13 ,\tt2_reg[15]_i_1_n_14 ,\tt2_reg[15]_i_1_n_15 }),
        .S({\tt2[15]_i_2_n_0 ,\tt2[15]_i_3_n_0 ,\tt2[15]_i_4_n_0 ,\tt2[15]_i_5_n_0 ,\tt2[15]_i_6_n_0 ,\tt2[15]_i_7_n_0 ,\tt2[15]_i_8_n_0 ,\tt2[15]_i_9_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[16] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[20]_i_1_n_15 ),
        .Q(tt2[16]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[17] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[20]_i_1_n_14 ),
        .Q(tt2[17]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[18] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[20]_i_1_n_13 ),
        .Q(tt2[18]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[19] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[20]_i_1_n_12 ),
        .Q(tt2[19]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[1] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_14 ),
        .Q(tt2[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[20] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[20]_i_1_n_11 ),
        .Q(tt2[20]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tt2_reg[20]_i_1 
       (.CI(\tt2_reg[15]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_tt2_reg[20]_i_1_CO_UNCONNECTED [7:4],\tt2_reg[20]_i_1_n_4 ,\tt2_reg[20]_i_1_n_5 ,\tt2_reg[20]_i_1_n_6 ,\tt2_reg[20]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,R[18],\tt2[20]_i_2_n_0 ,dd2__0[18],dd2__0[16]}),
        .O({\NLW_tt2_reg[20]_i_1_O_UNCONNECTED [7:5],\tt2_reg[20]_i_1_n_11 ,\tt2_reg[20]_i_1_n_12 ,\tt2_reg[20]_i_1_n_13 ,\tt2_reg[20]_i_1_n_14 ,\tt2_reg[20]_i_1_n_15 }),
        .S({1'b0,1'b0,1'b0,\tt2[20]_i_3_n_0 ,\tt2[20]_i_4_n_0 ,\tt2[20]_i_5_n_0 ,\tt2[20]_i_6_n_0 ,\tt2[20]_i_7_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[2] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_13 ),
        .Q(tt2[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[3] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_12 ),
        .Q(tt2[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[4] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_11 ),
        .Q(tt2[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[5] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_10 ),
        .Q(tt2[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[6] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_9 ),
        .Q(tt2[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[7] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[7]_i_1_n_8 ),
        .Q(tt2[7]),
        .R(1'b0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tt2_reg[7]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\tt2_reg[7]_i_1_n_0 ,\tt2_reg[7]_i_1_n_1 ,\tt2_reg[7]_i_1_n_2 ,\tt2_reg[7]_i_1_n_3 ,\tt2_reg[7]_i_1_n_4 ,\tt2_reg[7]_i_1_n_5 ,\tt2_reg[7]_i_1_n_6 ,\tt2_reg[7]_i_1_n_7 }),
        .DI(dd2[7:0]),
        .O({\tt2_reg[7]_i_1_n_8 ,\tt2_reg[7]_i_1_n_9 ,\tt2_reg[7]_i_1_n_10 ,\tt2_reg[7]_i_1_n_11 ,\tt2_reg[7]_i_1_n_12 ,\tt2_reg[7]_i_1_n_13 ,\tt2_reg[7]_i_1_n_14 ,\tt2_reg[7]_i_1_n_15 }),
        .S({\tt2[7]_i_2_n_0 ,\tt2[7]_i_3_n_0 ,\tt2[7]_i_4_n_0 ,\tt2[7]_i_5_n_0 ,\tt2[7]_i_6_n_0 ,\tt2[7]_i_7_n_0 ,\tt2[7]_i_8_n_0 ,\tt2[7]_i_9_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[8] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_15 ),
        .Q(tt2[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tt2_reg[9] 
       (.C(clk_i),
        .CE(E),
        .D(\tt2_reg[15]_i_1_n_14 ),
        .Q(tt2[9]),
        .R(1'b0));
  LUT1 #(
    .INIT(2'h1)) 
    \tt2_z1[21]_i_2 
       (.I0(tt2[20]),
        .O(\tt2_z1[21]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \tt2_z1[21]_i_3 
       (.I0(tt2[19]),
        .O(\tt2_z1[21]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \tt2_z1[21]_i_4 
       (.I0(tt2[18]),
        .O(\tt2_z1[21]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \tt2_z1[21]_i_5 
       (.I0(tt2[17]),
        .O(\tt2_z1[21]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \tt2_z1[21]_i_6 
       (.I0(tt2[16]),
        .O(\tt2_z1[21]_i_6_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_27),
        .Q(tt2_z1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_26),
        .Q(tt2_z1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_25),
        .Q(tt2_z1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_24),
        .Q(tt2_z1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_23),
        .Q(tt2_z1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_22),
        .Q(tt2_z1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_21),
        .Q(tt2_z1[16]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_20),
        .Q(tt2_z1[17]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_19),
        .Q(tt2_z1[18]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_18),
        .Q(tt2_z1[19]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_17),
        .Q(tt2_z1[20]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_16),
        .Q(tt2_z1[21]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_33),
        .Q(tt2_z1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_32),
        .Q(tt2_z1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_31),
        .Q(tt2_z1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_30),
        .Q(tt2_z1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_29),
        .Q(tt2_z1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2_z1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(DZ1_n_28),
        .Q(tt2_z1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[0]),
        .Q(tt2d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[10]),
        .Q(tt2d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[11]),
        .Q(tt2d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[12]),
        .Q(tt2d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[13]),
        .Q(tt2d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[14]),
        .Q(tt2d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[15]),
        .Q(tt2d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[1]),
        .Q(tt2d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[2]),
        .Q(tt2d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[3]),
        .Q(tt2d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[4]),
        .Q(tt2d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[5]),
        .Q(tt2d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[6]),
        .Q(tt2d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[7]),
        .Q(tt2d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[8]),
        .Q(tt2d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2[9]),
        .Q(tt2d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[0]),
        .Q(tt2d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[10]),
        .Q(tt2d2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[11]),
        .Q(tt2d2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[12]),
        .Q(tt2d2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[13]),
        .Q(tt2d2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[14]),
        .Q(tt2d2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[15]),
        .Q(tt2d2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[1]),
        .Q(tt2d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[2]),
        .Q(tt2d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[3]),
        .Q(tt2d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[4]),
        .Q(tt2d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[5]),
        .Q(tt2d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[6]),
        .Q(tt2d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[7]),
        .Q(tt2d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[8]),
        .Q(tt2d2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \tt2d2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(tt2d1[9]),
        .Q(tt2d2[9]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[0]),
        .Q(z1d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[10]),
        .Q(z1d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[11]),
        .Q(z1d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[12]),
        .Q(z1d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[13]),
        .Q(z1d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[14]),
        .Q(z1d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[15]),
        .Q(z1d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[1]),
        .Q(z1d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[2]),
        .Q(z1d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[3]),
        .Q(z1d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[4]),
        .Q(z1d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[5]),
        .Q(z1d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[6]),
        .Q(z1d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[7]),
        .Q(z1d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[8]),
        .Q(z1d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1[9]),
        .Q(z1d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[0]),
        .Q(z1d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[10]),
        .Q(z1d2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[11]),
        .Q(z1d2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[12]),
        .Q(z1d2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[13]),
        .Q(z1d2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[14]),
        .Q(z1d2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[15]),
        .Q(z1d2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[1]),
        .Q(z1d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[2]),
        .Q(z1d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[3]),
        .Q(z1d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[4]),
        .Q(z1d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[5]),
        .Q(z1d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[6]),
        .Q(z1d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[7]),
        .Q(z1d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[8]),
        .Q(z1d2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \z1d2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z1d1[9]),
        .Q(z1d2[9]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[0]),
        .Q(z2d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[10]),
        .Q(z2d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[11]),
        .Q(z2d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[12]),
        .Q(z2d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[13]),
        .Q(z2d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[14]),
        .Q(z2d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[15]),
        .Q(z2d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[1]),
        .Q(z2d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[2]),
        .Q(z2d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[3]),
        .Q(z2d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[4]),
        .Q(z2d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[5]),
        .Q(z2d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[6]),
        .Q(z2d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[7]),
        .Q(z2d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[8]),
        .Q(z2d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2[9]),
        .Q(z2d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[0]),
        .Q(z2d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[10]),
        .Q(z2d2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[11]),
        .Q(z2d2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[12]),
        .Q(z2d2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[13]),
        .Q(z2d2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[14]),
        .Q(z2d2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[15]),
        .Q(z2d2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[1]),
        .Q(z2d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[2]),
        .Q(z2d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[3]),
        .Q(z2d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[4]),
        .Q(z2d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[5]),
        .Q(z2d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[6]),
        .Q(z2d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[7]),
        .Q(z2d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[8]),
        .Q(z2d2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \z2d2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z2d1[9]),
        .Q(z2d2[9]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[0]),
        .Q(z3d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[10]),
        .Q(z3d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[11]),
        .Q(z3d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[12]),
        .Q(z3d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[13]),
        .Q(z3d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[14]),
        .Q(z3d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[15]),
        .Q(z3d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[1]),
        .Q(z3d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[2]),
        .Q(z3d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[3]),
        .Q(z3d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[4]),
        .Q(z3d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[5]),
        .Q(z3d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[6]),
        .Q(z3d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[7]),
        .Q(z3d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[8]),
        .Q(z3d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3[9]),
        .Q(z3d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[0]),
        .Q(z3d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[10]),
        .Q(z3d2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[11]),
        .Q(z3d2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[12]),
        .Q(z3d2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[13]),
        .Q(z3d2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[14]),
        .Q(z3d2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[15]),
        .Q(z3d2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[1]),
        .Q(z3d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[2]),
        .Q(z3d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[3]),
        .Q(z3d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[4]),
        .Q(z3d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[5]),
        .Q(z3d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[6]),
        .Q(z3d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[7]),
        .Q(z3d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[8]),
        .Q(z3d2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \z3d2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(z3d1[9]),
        .Q(z3d2[9]));
endmodule

(* ORIG_REF_NAME = "SwitchAsyncFIFO" *) 
module switch_elements_SwitchAsyncFIFO
   (rst_i_0,
    this_cycle,
    D,
    E,
    \qvDataOut_reg[71] ,
    \qvDataOut_reg[69] ,
    \qvDataOut_reg[62] ,
    get_sfd0,
    \qvDataOut_reg[45] ,
    clk_i,
    Q,
    rst_i,
    recv_rst,
    MemDataIn);
  output rst_i_0;
  output this_cycle;
  output [5:0]D;
  output [0:0]E;
  output [71:0]\qvDataOut_reg[71] ;
  output [2:0]\qvDataOut_reg[69] ;
  output [7:0]\qvDataOut_reg[62] ;
  output get_sfd0;
  output \qvDataOut_reg[45] ;
  input clk_i;
  input [0:0]Q;
  input rst_i;
  input recv_rst;
  input [71:0]MemDataIn;

  wire [5:0]D;
  wire [0:0]E;
  wire [71:0]MemDataIn;
  wire [71:0]MemDataOut;
  wire MemWEn;
  wire [0:0]Q;
  wire clk_i;
  wire get_sfd0;
  wire \qvDataOut_reg[45] ;
  wire [7:0]\qvDataOut_reg[62] ;
  wire [2:0]\qvDataOut_reg[69] ;
  wire [71:0]\qvDataOut_reg[71] ;
  wire recv_rst;
  wire rst_i;
  wire rst_i_0;
  wire this_cycle;
  wire [4:0]vReadAddr;
  wire [4:0]vWAddr;

  switch_elements_FifoControl_ASYN Fifo_Controller
       (.ADDRH(vWAddr),
        .D(vReadAddr),
        .E(MemWEn),
        .Q(Q),
        .clk_i(clk_i),
        .get_sfd0(get_sfd0),
        .\qvDataOut_reg[25]_0 (D),
        .\qvDataOut_reg[45]_0 (\qvDataOut_reg[45] ),
        .\qvDataOut_reg[62]_0 (\qvDataOut_reg[62] ),
        .\qvDataOut_reg[66]_0 (E),
        .\qvDataOut_reg[69]_0 (\qvDataOut_reg[69] ),
        .\qvDataOut_reg[71]_0 (\qvDataOut_reg[71] ),
        .\qvDataOut_reg[71]_1 (MemDataOut),
        .recv_rst(recv_rst),
        .rst_i(rst_i),
        .rst_i_0(rst_i_0),
        .this_cycle(this_cycle));
  switch_elements_DualPortRAM_ASYN Fifo_Storage
       (.ADDRH(vWAddr),
        .D(vReadAddr),
        .E(MemWEn),
        .MemDataIn(MemDataIn),
        .clk_i(clk_i),
        .clk_i_0(MemDataOut));
endmodule

(* ORIG_REF_NAME = "SwitchSyncFIFO" *) 
module switch_elements_SwitchSyncFIFO
   (rxfifo_empty,
    D,
    pad_cnt_reg1,
    fifo_rd_en,
    qEmpty_reg,
    \ovDataOut_reg[63]_0 ,
    \qvRAddr_reg[6] ,
    receiving_d2,
    Q,
    \pad_cnt_reg_reg[0] ,
    fifo_rd_en_reg,
    \pad_rxc_reg_reg[0] ,
    fifo_rd_en_reg_0,
    pad_frame_d1_reg,
    clk_i,
    rxd64_d3,
    reset_dcm);
  output rxfifo_empty;
  output [2:0]D;
  output pad_cnt_reg1;
  output fifo_rd_en;
  output qEmpty_reg;
  output [63:0]\ovDataOut_reg[63]_0 ;
  input \qvRAddr_reg[6] ;
  input receiving_d2;
  input [2:0]Q;
  input [2:0]\pad_cnt_reg_reg[0] ;
  input [1:0]fifo_rd_en_reg;
  input \pad_rxc_reg_reg[0] ;
  input fifo_rd_en_reg_0;
  input pad_frame_d1_reg;
  input clk_i;
  input [63:0]rxd64_d3;
  input reset_dcm;

  wire [2:0]D;
  wire Fifo_Ctrl_n_10;
  wire Fifo_Ctrl_n_11;
  wire Fifo_Ctrl_n_20;
  wire Fifo_Ctrl_n_21;
  wire Fifo_Ctrl_n_5;
  wire Fifo_Ctrl_n_6;
  wire Fifo_Ctrl_n_7;
  wire Fifo_Ctrl_n_8;
  wire Fifo_Ctrl_n_9;
  wire [2:0]Q;
  wire clk_i;
  wire fifo_rd_en;
  wire [1:0]fifo_rd_en_reg;
  wire fifo_rd_en_reg_0;
  wire \ovDataOut[63]_i_1_n_0 ;
  wire [63:0]ovDataOut_i;
  wire [63:0]\ovDataOut_reg[63]_0 ;
  wire pad_cnt_reg1;
  wire [2:0]\pad_cnt_reg_reg[0] ;
  wire pad_frame_d1_reg;
  wire \pad_rxc_reg_reg[0] ;
  wire qEmpty_reg;
  wire \qvRAddr_reg[6] ;
  wire [5:0]qvWAddr;
  wire receiving_d2;
  wire reset_dcm;
  wire [63:0]rxd64_d3;
  wire rxfifo_empty;

  switch_elements_FifoControl Fifo_Ctrl
       (.D(D),
        .\FSM_sequential_fifo_state_reg[0] (pad_cnt_reg1),
        .Q(Q),
        .clk_i(clk_i),
        .fifo_rd_en(fifo_rd_en),
        .fifo_rd_en_reg(fifo_rd_en_reg),
        .fifo_rd_en_reg_0(fifo_rd_en_reg_0),
        .\pad_cnt_reg_reg[0] (\pad_cnt_reg_reg[0] ),
        .pad_frame_d1_reg(pad_frame_d1_reg),
        .\pad_rxc_reg_reg[0] (\pad_rxc_reg_reg[0] ),
        .qEmpty_reg_0(rxfifo_empty),
        .qEmpty_reg_1(qEmpty_reg),
        .qFull_reg_0(Fifo_Ctrl_n_20),
        .qFull_reg_1(Fifo_Ctrl_n_21),
        .\qvRAddr_reg[6]_0 ({Fifo_Ctrl_n_5,Fifo_Ctrl_n_6,Fifo_Ctrl_n_7,Fifo_Ctrl_n_8,Fifo_Ctrl_n_9,Fifo_Ctrl_n_10,Fifo_Ctrl_n_11}),
        .\qvRAddr_reg[6]_1 (\qvRAddr_reg[6] ),
        .\qvWAddr_reg[5]_0 (qvWAddr),
        .receiving_d2(receiving_d2),
        .reset_dcm(reset_dcm));
  switch_elements_DualPortRAM Fifo_Storage
       (.clk_i(clk_i),
        .ovDataOut_i(ovDataOut_i),
        .\ovDataOut_reg[0] ({Fifo_Ctrl_n_5,Fifo_Ctrl_n_6,Fifo_Ctrl_n_7,Fifo_Ctrl_n_8,Fifo_Ctrl_n_9,Fifo_Ctrl_n_10,Fifo_Ctrl_n_11}),
        .\ovDataOut_reg[0]_0 (Fifo_Ctrl_n_21),
        .\ovDataOut_reg[63] (qvWAddr),
        .\ovDataOut_reg[63]_0 (Fifo_Ctrl_n_20),
        .rxd64_d3(rxd64_d3));
  LUT2 #(
    .INIT(4'hB)) 
    \ovDataOut[63]_i_1 
       (.I0(rxfifo_empty),
        .I1(\qvRAddr_reg[6] ),
        .O(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[0]),
        .Q(\ovDataOut_reg[63]_0 [0]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[10]),
        .Q(\ovDataOut_reg[63]_0 [10]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[11]),
        .Q(\ovDataOut_reg[63]_0 [11]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[12]),
        .Q(\ovDataOut_reg[63]_0 [12]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[13]),
        .Q(\ovDataOut_reg[63]_0 [13]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[14]),
        .Q(\ovDataOut_reg[63]_0 [14]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[15]),
        .Q(\ovDataOut_reg[63]_0 [15]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[16]),
        .Q(\ovDataOut_reg[63]_0 [16]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[17]),
        .Q(\ovDataOut_reg[63]_0 [17]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[18]),
        .Q(\ovDataOut_reg[63]_0 [18]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[19]),
        .Q(\ovDataOut_reg[63]_0 [19]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[1]),
        .Q(\ovDataOut_reg[63]_0 [1]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[20]),
        .Q(\ovDataOut_reg[63]_0 [20]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[21]),
        .Q(\ovDataOut_reg[63]_0 [21]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[22]),
        .Q(\ovDataOut_reg[63]_0 [22]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[23]),
        .Q(\ovDataOut_reg[63]_0 [23]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[24]),
        .Q(\ovDataOut_reg[63]_0 [24]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[25]),
        .Q(\ovDataOut_reg[63]_0 [25]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[26]),
        .Q(\ovDataOut_reg[63]_0 [26]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[27]),
        .Q(\ovDataOut_reg[63]_0 [27]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[28]),
        .Q(\ovDataOut_reg[63]_0 [28]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[29]),
        .Q(\ovDataOut_reg[63]_0 [29]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[2]),
        .Q(\ovDataOut_reg[63]_0 [2]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[30]),
        .Q(\ovDataOut_reg[63]_0 [30]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[31]),
        .Q(\ovDataOut_reg[63]_0 [31]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[32]),
        .Q(\ovDataOut_reg[63]_0 [32]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[33]),
        .Q(\ovDataOut_reg[63]_0 [33]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[34]),
        .Q(\ovDataOut_reg[63]_0 [34]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[35]),
        .Q(\ovDataOut_reg[63]_0 [35]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[36]),
        .Q(\ovDataOut_reg[63]_0 [36]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[37]),
        .Q(\ovDataOut_reg[63]_0 [37]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[38]),
        .Q(\ovDataOut_reg[63]_0 [38]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[39]),
        .Q(\ovDataOut_reg[63]_0 [39]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[3]),
        .Q(\ovDataOut_reg[63]_0 [3]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[40]),
        .Q(\ovDataOut_reg[63]_0 [40]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[41]),
        .Q(\ovDataOut_reg[63]_0 [41]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[42]),
        .Q(\ovDataOut_reg[63]_0 [42]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[43]),
        .Q(\ovDataOut_reg[63]_0 [43]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[44]),
        .Q(\ovDataOut_reg[63]_0 [44]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[45]),
        .Q(\ovDataOut_reg[63]_0 [45]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[46]),
        .Q(\ovDataOut_reg[63]_0 [46]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[47]),
        .Q(\ovDataOut_reg[63]_0 [47]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[48]),
        .Q(\ovDataOut_reg[63]_0 [48]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[49]),
        .Q(\ovDataOut_reg[63]_0 [49]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[4]),
        .Q(\ovDataOut_reg[63]_0 [4]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[50]),
        .Q(\ovDataOut_reg[63]_0 [50]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[51]),
        .Q(\ovDataOut_reg[63]_0 [51]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[52]),
        .Q(\ovDataOut_reg[63]_0 [52]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[53]),
        .Q(\ovDataOut_reg[63]_0 [53]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[54]),
        .Q(\ovDataOut_reg[63]_0 [54]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[55]),
        .Q(\ovDataOut_reg[63]_0 [55]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[56]),
        .Q(\ovDataOut_reg[63]_0 [56]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[57]),
        .Q(\ovDataOut_reg[63]_0 [57]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[58]),
        .Q(\ovDataOut_reg[63]_0 [58]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[59]),
        .Q(\ovDataOut_reg[63]_0 [59]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[5]),
        .Q(\ovDataOut_reg[63]_0 [5]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[60]),
        .Q(\ovDataOut_reg[63]_0 [60]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[61]),
        .Q(\ovDataOut_reg[63]_0 [61]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[62]),
        .Q(\ovDataOut_reg[63]_0 [62]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[63]),
        .Q(\ovDataOut_reg[63]_0 [63]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[6]),
        .Q(\ovDataOut_reg[63]_0 [6]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[7]),
        .Q(\ovDataOut_reg[63]_0 [7]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[8]),
        .Q(\ovDataOut_reg[63]_0 [8]),
        .R(\ovDataOut[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[9]),
        .Q(\ovDataOut_reg[63]_0 [9]),
        .R(\ovDataOut[63]_i_1_n_0 ));
endmodule

(* ORIG_REF_NAME = "SwitchSyncFIFO" *) 
module switch_elements_SwitchSyncFIFO__parameterized0
   (D,
    \ovDataOut_reg[5]_0 ,
    \ovDataOut_reg[7]_0 ,
    \qvRAddr_reg[6] ,
    receiving_d2,
    rxfifo_empty,
    Q,
    bad_frame_get,
    good_frame_get,
    \rx_data_valid_reg[1] ,
    \rx_data_valid_reg[7] ,
    \rx_data_valid_reg[6] ,
    \rx_data_valid_reg[1]_0 ,
    \rx_data_valid_reg[7]_0 ,
    \rx_data_valid_reg[0] ,
    clk_i,
    vDataIn,
    reset_dcm);
  output [1:0]D;
  output \ovDataOut_reg[5]_0 ;
  output [7:0]\ovDataOut_reg[7]_0 ;
  input \qvRAddr_reg[6] ;
  input receiving_d2;
  input rxfifo_empty;
  input [1:0]Q;
  input bad_frame_get;
  input good_frame_get;
  input \rx_data_valid_reg[1] ;
  input [2:0]\rx_data_valid_reg[7] ;
  input [6:0]\rx_data_valid_reg[6] ;
  input \rx_data_valid_reg[1]_0 ;
  input \rx_data_valid_reg[7]_0 ;
  input \rx_data_valid_reg[0] ;
  input clk_i;
  input [7:0]vDataIn;
  input reset_dcm;

  wire [1:0]D;
  wire \FSM_sequential_fifo_state[1]_i_4_n_0 ;
  wire Fifo_Ctrl_n_0;
  wire Fifo_Ctrl_n_1;
  wire Fifo_Ctrl_n_10;
  wire Fifo_Ctrl_n_11;
  wire Fifo_Ctrl_n_12;
  wire Fifo_Ctrl_n_13;
  wire Fifo_Ctrl_n_14;
  wire Fifo_Ctrl_n_15;
  wire Fifo_Ctrl_n_2;
  wire Fifo_Ctrl_n_3;
  wire Fifo_Ctrl_n_4;
  wire Fifo_Ctrl_n_5;
  wire Fifo_Ctrl_n_6;
  wire Fifo_Ctrl_n_7;
  wire Fifo_Ctrl_n_8;
  wire Fifo_Ctrl_n_9;
  wire [1:0]Q;
  wire bad_frame_get;
  wire clk_i;
  wire good_frame_get;
  wire \ovDataOut[7]_i_1_n_0 ;
  wire [7:0]ovDataOut_i;
  wire \ovDataOut_reg[5]_0 ;
  wire [7:0]\ovDataOut_reg[7]_0 ;
  wire \qvRAddr_reg[6] ;
  wire receiving_d2;
  wire reset_dcm;
  wire \rx_data_valid_reg[0] ;
  wire \rx_data_valid_reg[1] ;
  wire \rx_data_valid_reg[1]_0 ;
  wire [6:0]\rx_data_valid_reg[6] ;
  wire [2:0]\rx_data_valid_reg[7] ;
  wire \rx_data_valid_reg[7]_0 ;
  wire [7:0]rx_data_valid_tmp;
  wire rxfifo_empty;
  wire [7:0]vDataIn;

  LUT6 #(
    .INIT(64'h5F5F5F5D57575755)) 
    \FSM_sequential_fifo_state[0]_i_1 
       (.I0(\ovDataOut_reg[5]_0 ),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(bad_frame_get),
        .I4(good_frame_get),
        .I5(rxfifo_empty),
        .O(D[0]));
  LUT4 #(
    .INIT(16'h5F75)) 
    \FSM_sequential_fifo_state[1]_i_1 
       (.I0(\ovDataOut_reg[5]_0 ),
        .I1(rxfifo_empty),
        .I2(Q[0]),
        .I3(Q[1]),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \FSM_sequential_fifo_state[1]_i_3 
       (.I0(\FSM_sequential_fifo_state[1]_i_4_n_0 ),
        .I1(rx_data_valid_tmp[5]),
        .I2(rx_data_valid_tmp[4]),
        .I3(rx_data_valid_tmp[6]),
        .I4(rx_data_valid_tmp[7]),
        .I5(Q[1]),
        .O(\ovDataOut_reg[5]_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \FSM_sequential_fifo_state[1]_i_4 
       (.I0(rx_data_valid_tmp[1]),
        .I1(rx_data_valid_tmp[0]),
        .I2(rx_data_valid_tmp[3]),
        .I3(rx_data_valid_tmp[2]),
        .O(\FSM_sequential_fifo_state[1]_i_4_n_0 ));
  switch_elements_FifoControl_2 Fifo_Ctrl
       (.Q({Fifo_Ctrl_n_1,Fifo_Ctrl_n_2,Fifo_Ctrl_n_3,Fifo_Ctrl_n_4,Fifo_Ctrl_n_5,Fifo_Ctrl_n_6,Fifo_Ctrl_n_7}),
        .clk_i(clk_i),
        .qEmpty_reg_0(Fifo_Ctrl_n_0),
        .qFull_reg_0(Fifo_Ctrl_n_14),
        .qFull_reg_1(Fifo_Ctrl_n_15),
        .\qvRAddr_reg[6]_0 (\qvRAddr_reg[6] ),
        .\qvWAddr_reg[5]_0 ({Fifo_Ctrl_n_8,Fifo_Ctrl_n_9,Fifo_Ctrl_n_10,Fifo_Ctrl_n_11,Fifo_Ctrl_n_12,Fifo_Ctrl_n_13}),
        .receiving_d2(receiving_d2),
        .reset_dcm(reset_dcm));
  switch_elements_DualPortRAM__parameterized0 Fifo_Storage
       (.Q({Fifo_Ctrl_n_1,Fifo_Ctrl_n_2,Fifo_Ctrl_n_3,Fifo_Ctrl_n_4,Fifo_Ctrl_n_5,Fifo_Ctrl_n_6,Fifo_Ctrl_n_7}),
        .clk_i(clk_i),
        .ovDataOut_i(ovDataOut_i),
        .\ovDataOut_reg[0] (Fifo_Ctrl_n_14),
        .\ovDataOut_reg[7] ({Fifo_Ctrl_n_8,Fifo_Ctrl_n_9,Fifo_Ctrl_n_10,Fifo_Ctrl_n_11,Fifo_Ctrl_n_12,Fifo_Ctrl_n_13}),
        .\ovDataOut_reg[7]_0 (Fifo_Ctrl_n_15),
        .vDataIn(vDataIn));
  LUT2 #(
    .INIT(4'hB)) 
    \ovDataOut[7]_i_1 
       (.I0(Fifo_Ctrl_n_0),
        .I1(\qvRAddr_reg[6] ),
        .O(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[0]),
        .Q(rx_data_valid_tmp[0]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[1]),
        .Q(rx_data_valid_tmp[1]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[2]),
        .Q(rx_data_valid_tmp[2]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[3]),
        .Q(rx_data_valid_tmp[3]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[4]),
        .Q(rx_data_valid_tmp[4]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[5]),
        .Q(rx_data_valid_tmp[5]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[6]),
        .Q(rx_data_valid_tmp[6]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \ovDataOut_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(ovDataOut_i[7]),
        .Q(rx_data_valid_tmp[7]),
        .R(\ovDataOut[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8F800000FF000000)) 
    \rx_data_valid[0]_i_1 
       (.I0(\rx_data_valid_reg[7] [0]),
        .I1(\rx_data_valid_reg[6] [0]),
        .I2(\rx_data_valid_reg[0] ),
        .I3(rx_data_valid_tmp[0]),
        .I4(Q[1]),
        .I5(\rx_data_valid_reg[7]_0 ),
        .O(\ovDataOut_reg[7]_0 [0]));
  LUT5 #(
    .INIT(32'hF4444444)) 
    \rx_data_valid[1]_i_1 
       (.I0(\rx_data_valid_reg[1] ),
        .I1(rx_data_valid_tmp[1]),
        .I2(\rx_data_valid_reg[7] [0]),
        .I3(\rx_data_valid_reg[6] [1]),
        .I4(\rx_data_valid_reg[1]_0 ),
        .O(\ovDataOut_reg[7]_0 [1]));
  LUT5 #(
    .INIT(32'hF4444444)) 
    \rx_data_valid[2]_i_1 
       (.I0(\rx_data_valid_reg[1] ),
        .I1(rx_data_valid_tmp[2]),
        .I2(\rx_data_valid_reg[7] [0]),
        .I3(\rx_data_valid_reg[6] [2]),
        .I4(\rx_data_valid_reg[1]_0 ),
        .O(\ovDataOut_reg[7]_0 [2]));
  LUT5 #(
    .INIT(32'hF4444444)) 
    \rx_data_valid[3]_i_1 
       (.I0(\rx_data_valid_reg[1] ),
        .I1(rx_data_valid_tmp[3]),
        .I2(\rx_data_valid_reg[7] [0]),
        .I3(\rx_data_valid_reg[6] [3]),
        .I4(\rx_data_valid_reg[1]_0 ),
        .O(\ovDataOut_reg[7]_0 [3]));
  LUT5 #(
    .INIT(32'hF4444444)) 
    \rx_data_valid[4]_i_1 
       (.I0(\rx_data_valid_reg[1] ),
        .I1(rx_data_valid_tmp[4]),
        .I2(\rx_data_valid_reg[7] [0]),
        .I3(\rx_data_valid_reg[6] [4]),
        .I4(\rx_data_valid_reg[1]_0 ),
        .O(\ovDataOut_reg[7]_0 [4]));
  LUT5 #(
    .INIT(32'hF4444444)) 
    \rx_data_valid[5]_i_1 
       (.I0(\rx_data_valid_reg[1] ),
        .I1(rx_data_valid_tmp[5]),
        .I2(\rx_data_valid_reg[7] [0]),
        .I3(\rx_data_valid_reg[6] [5]),
        .I4(\rx_data_valid_reg[1]_0 ),
        .O(\ovDataOut_reg[7]_0 [5]));
  LUT5 #(
    .INIT(32'hF4444444)) 
    \rx_data_valid[6]_i_1 
       (.I0(\rx_data_valid_reg[1] ),
        .I1(rx_data_valid_tmp[6]),
        .I2(\rx_data_valid_reg[7] [0]),
        .I3(\rx_data_valid_reg[6] [6]),
        .I4(\rx_data_valid_reg[1]_0 ),
        .O(\ovDataOut_reg[7]_0 [6]));
  LUT5 #(
    .INIT(32'h88888808)) 
    \rx_data_valid[7]_i_1 
       (.I0(rx_data_valid_tmp[7]),
        .I1(Q[1]),
        .I2(\rx_data_valid_reg[7]_0 ),
        .I3(\rx_data_valid_reg[7] [2]),
        .I4(\rx_data_valid_reg[7] [1]),
        .O(\ovDataOut_reg[7]_0 [7]));
endmodule

(* ORIG_REF_NAME = "TRANSMIT_TOP" *) 
module switch_elements_TRANSMIT_TOP
   (E,
    TX_ACK,
    TX_STATS_VALID,
    TXSTATREGPLUS,
    TXD,
    TXC,
    FC_TRANS_PAUSEVAL,
    clk_i,
    rst_i,
    out,
    load_final_CRC_reg_0,
    TX_CFG_REG_VALID,
    TX_CFG_REG_VALUE,
    FC_TRANS_PAUSEDATA,
    TX_DATA,
    \TX_DATA_VALID_REG_reg[7]_0 ,
    apply_pause_delay_reg_0,
    tx_undderrun_int_reg_0,
    I94,
    \DELAY_ACK_reg[7]_0 );
  output [0:0]E;
  output TX_ACK;
  output TX_STATS_VALID;
  output [24:0]TXSTATREGPLUS;
  output [63:0]TXD;
  output [7:0]TXC;
  input FC_TRANS_PAUSEVAL;
  input clk_i;
  input rst_i;
  input out;
  input load_final_CRC_reg_0;
  input TX_CFG_REG_VALID;
  input [3:0]TX_CFG_REG_VALUE;
  input [15:0]FC_TRANS_PAUSEDATA;
  input [63:0]TX_DATA;
  input [7:0]\TX_DATA_VALID_REG_reg[7]_0 ;
  input apply_pause_delay_reg_0;
  input tx_undderrun_int_reg_0;
  input [15:0]I94;
  input [7:0]\DELAY_ACK_reg[7]_0 ;

  wire [15:2]BYTE_COUNTER;
  wire [31:0]CRC_32_64;
  wire [15:0]DELAY_ACK;
  wire \DELAY_ACK[0]_i_1_n_0 ;
  wire \DELAY_ACK[10]_i_1_n_0 ;
  wire \DELAY_ACK[11]_i_1_n_0 ;
  wire \DELAY_ACK[12]_i_1_n_0 ;
  wire \DELAY_ACK[13]_i_1_n_0 ;
  wire \DELAY_ACK[14]_i_1_n_0 ;
  wire \DELAY_ACK[15]_i_1_n_0 ;
  wire \DELAY_ACK[15]_i_2_n_0 ;
  wire \DELAY_ACK[1]_i_1_n_0 ;
  wire \DELAY_ACK[2]_i_1_n_0 ;
  wire \DELAY_ACK[3]_i_1_n_0 ;
  wire \DELAY_ACK[4]_i_1_n_0 ;
  wire \DELAY_ACK[5]_i_1_n_0 ;
  wire \DELAY_ACK[6]_i_1_n_0 ;
  wire \DELAY_ACK[7]_i_1_n_0 ;
  wire \DELAY_ACK[8]_i_1_n_0 ;
  wire \DELAY_ACK[9]_i_1_n_0 ;
  wire [7:0]\DELAY_ACK_reg[7]_0 ;
  wire [0:0]E;
  wire [15:0]FC_TRANS_PAUSEDATA;
  wire FC_TRANS_PAUSEVAL;
  wire FRAME_START;
  wire FRAME_START_i_3_n_0;
  wire FRAME_START_i_4_n_0;
  wire [15:0]I94;
  wire [4:2]MAX_FRAME_SIZE;
  wire \MAX_FRAME_SIZE[2]_i_1_n_0 ;
  wire \MAX_FRAME_SIZE[3]_i_1_n_0 ;
  wire \MAX_FRAME_SIZE[4]_i_1_n_0 ;
  wire \OVERFLOW_DATA[17]_i_2_n_0 ;
  wire \OVERFLOW_DATA[23]_i_2_n_0 ;
  wire \OVERFLOW_DATA[25]_i_1_n_0 ;
  wire \OVERFLOW_DATA[31]_i_1_n_0 ;
  wire \OVERFLOW_DATA[31]_i_2_n_0 ;
  wire \OVERFLOW_DATA[33]_i_1_n_0 ;
  wire \OVERFLOW_DATA[39]_i_1_n_0 ;
  wire \OVERFLOW_DATA[39]_i_2_n_0 ;
  wire \OVERFLOW_DATA[8]_i_2_n_0 ;
  wire \OVERFLOW_DATA_reg_n_0_[0] ;
  wire \OVERFLOW_DATA_reg_n_0_[10] ;
  wire \OVERFLOW_DATA_reg_n_0_[11] ;
  wire \OVERFLOW_DATA_reg_n_0_[12] ;
  wire \OVERFLOW_DATA_reg_n_0_[13] ;
  wire \OVERFLOW_DATA_reg_n_0_[14] ;
  wire \OVERFLOW_DATA_reg_n_0_[15] ;
  wire \OVERFLOW_DATA_reg_n_0_[16] ;
  wire \OVERFLOW_DATA_reg_n_0_[17] ;
  wire \OVERFLOW_DATA_reg_n_0_[18] ;
  wire \OVERFLOW_DATA_reg_n_0_[19] ;
  wire \OVERFLOW_DATA_reg_n_0_[1] ;
  wire \OVERFLOW_DATA_reg_n_0_[20] ;
  wire \OVERFLOW_DATA_reg_n_0_[21] ;
  wire \OVERFLOW_DATA_reg_n_0_[22] ;
  wire \OVERFLOW_DATA_reg_n_0_[23] ;
  wire \OVERFLOW_DATA_reg_n_0_[25] ;
  wire \OVERFLOW_DATA_reg_n_0_[2] ;
  wire \OVERFLOW_DATA_reg_n_0_[31] ;
  wire \OVERFLOW_DATA_reg_n_0_[33] ;
  wire \OVERFLOW_DATA_reg_n_0_[39] ;
  wire \OVERFLOW_DATA_reg_n_0_[3] ;
  wire \OVERFLOW_DATA_reg_n_0_[4] ;
  wire \OVERFLOW_DATA_reg_n_0_[5] ;
  wire \OVERFLOW_DATA_reg_n_0_[6] ;
  wire \OVERFLOW_DATA_reg_n_0_[7] ;
  wire \OVERFLOW_DATA_reg_n_0_[8] ;
  wire \OVERFLOW_DATA_reg_n_0_[9] ;
  wire \OVERFLOW_VALID[0]_i_1_n_0 ;
  wire \OVERFLOW_VALID[1]_i_1_n_0 ;
  wire \OVERFLOW_VALID[2]_i_1_n_0 ;
  wire \OVERFLOW_VALID[2]_i_2_n_0 ;
  wire \OVERFLOW_VALID[2]_i_3_n_0 ;
  wire [2:0]OVERFLOW_VALID__0;
  wire PAUSEVAL_DEL1_reg_srl2_n_0;
  wire PAUSEVAL_DEL2;
  wire RESET0;
  wire RESET02_out;
  wire [7:0]TXC;
  wire [63:0]TXD;
  wire [60:60]TXD_PAUSE_DEL1;
  wire [15:0]TXD_PAUSE_DEL2;
  wire [24:0]TXSTATREGPLUS;
  wire TX_ACK;
  wire TX_CFG_REG_VALID;
  wire [3:0]TX_CFG_REG_VALUE;
  wire [63:0]TX_DATA;
  wire [63:0]TX_DATA_DEL1;
  wire \TX_DATA_DEL11_reg[0]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[10]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[11]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[12]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[13]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[14]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[15]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[16]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[17]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[18]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[19]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[1]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[20]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[21]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[22]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[23]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[24]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[25]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[26]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[27]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[28]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[29]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[2]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[30]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[31]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[32]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[33]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[34]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[35]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[36]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[37]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[38]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[39]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[3]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[40]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[41]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[42]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[43]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[44]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[45]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[46]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[47]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[48]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[49]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[4]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[50]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[51]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[52]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[53]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[54]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[55]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[56]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[57]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[58]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[59]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[5]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[60]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[61]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[62]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[63]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[6]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[7]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[8]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL11_reg[9]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_DEL12_reg[0]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[10]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[11]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[12]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[13]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[14]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[15]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[16]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[17]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[18]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[19]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[1]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[20]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[21]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[22]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[23]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[24]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[25]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[26]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[27]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[28]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[29]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[2]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[30]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[31]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[32]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[33]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[34]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[35]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[36]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[37]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[38]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[39]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[3]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[40]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[41]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[42]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[43]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[44]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[45]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[46]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[47]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[48]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[49]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[4]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[50]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[51]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[52]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[53]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[54]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[55]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[56]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[57]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[58]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[59]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[5]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[60]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[61]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[62]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[63]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[6]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[7]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[8]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_DEL12_reg[9]_activity_blocks_c_8_n_0 ;
  wire [63:0]TX_DATA_DEL13;
  wire \TX_DATA_DEL14[15]_i_2_n_0 ;
  wire \TX_DATA_DEL14[18]_i_4_n_0 ;
  wire \TX_DATA_DEL14[23]_i_2_n_0 ;
  wire \TX_DATA_DEL14[25]_i_4_n_0 ;
  wire \TX_DATA_DEL14[33]_i_4_n_0 ;
  wire \TX_DATA_DEL14[33]_i_6_n_0 ;
  wire \TX_DATA_DEL14[39]_i_3_n_0 ;
  wire \TX_DATA_DEL14[39]_i_5_n_0 ;
  wire \TX_DATA_DEL14[41]_i_5_n_0 ;
  wire \TX_DATA_DEL14[47]_i_3_n_0 ;
  wire \TX_DATA_DEL14[48]_i_5_n_0 ;
  wire \TX_DATA_DEL14[48]_i_6_n_0 ;
  wire \TX_DATA_DEL14[49]_i_5_n_0 ;
  wire \TX_DATA_DEL14[49]_i_6_n_0 ;
  wire \TX_DATA_DEL14[50]_i_3_n_0 ;
  wire \TX_DATA_DEL14[50]_i_5_n_0 ;
  wire \TX_DATA_DEL14[51]_i_5_n_0 ;
  wire \TX_DATA_DEL14[52]_i_3_n_0 ;
  wire \TX_DATA_DEL14[53]_i_3_n_0 ;
  wire \TX_DATA_DEL14[54]_i_5_n_0 ;
  wire \TX_DATA_DEL14[54]_i_6_n_0 ;
  wire \TX_DATA_DEL14[55]_i_3_n_0 ;
  wire \TX_DATA_DEL14[57]_i_6_n_0 ;
  wire \TX_DATA_DEL14[57]_i_7_n_0 ;
  wire \TX_DATA_DEL14[57]_i_8_n_0 ;
  wire \TX_DATA_DEL14[58]_i_3_n_0 ;
  wire \TX_DATA_DEL14[58]_i_5_n_0 ;
  wire \TX_DATA_DEL14[58]_i_6_n_0 ;
  wire \TX_DATA_DEL14[58]_i_7_n_0 ;
  wire \TX_DATA_DEL14[63]_i_4_n_0 ;
  wire \TX_DATA_DEL14[63]_i_5_n_0 ;
  wire \TX_DATA_DEL14[63]_i_7_n_0 ;
  wire \TX_DATA_DEL14[63]_i_8_n_0 ;
  wire \TX_DATA_DEL14_reg_n_0_[0] ;
  wire \TX_DATA_DEL14_reg_n_0_[10] ;
  wire \TX_DATA_DEL14_reg_n_0_[11] ;
  wire \TX_DATA_DEL14_reg_n_0_[12] ;
  wire \TX_DATA_DEL14_reg_n_0_[13] ;
  wire \TX_DATA_DEL14_reg_n_0_[14] ;
  wire \TX_DATA_DEL14_reg_n_0_[15] ;
  wire \TX_DATA_DEL14_reg_n_0_[16] ;
  wire \TX_DATA_DEL14_reg_n_0_[17] ;
  wire \TX_DATA_DEL14_reg_n_0_[18] ;
  wire \TX_DATA_DEL14_reg_n_0_[19] ;
  wire \TX_DATA_DEL14_reg_n_0_[1] ;
  wire \TX_DATA_DEL14_reg_n_0_[20] ;
  wire \TX_DATA_DEL14_reg_n_0_[21] ;
  wire \TX_DATA_DEL14_reg_n_0_[22] ;
  wire \TX_DATA_DEL14_reg_n_0_[23] ;
  wire \TX_DATA_DEL14_reg_n_0_[24] ;
  wire \TX_DATA_DEL14_reg_n_0_[25] ;
  wire \TX_DATA_DEL14_reg_n_0_[26] ;
  wire \TX_DATA_DEL14_reg_n_0_[27] ;
  wire \TX_DATA_DEL14_reg_n_0_[28] ;
  wire \TX_DATA_DEL14_reg_n_0_[29] ;
  wire \TX_DATA_DEL14_reg_n_0_[2] ;
  wire \TX_DATA_DEL14_reg_n_0_[30] ;
  wire \TX_DATA_DEL14_reg_n_0_[31] ;
  wire \TX_DATA_DEL14_reg_n_0_[32] ;
  wire \TX_DATA_DEL14_reg_n_0_[33] ;
  wire \TX_DATA_DEL14_reg_n_0_[34] ;
  wire \TX_DATA_DEL14_reg_n_0_[35] ;
  wire \TX_DATA_DEL14_reg_n_0_[36] ;
  wire \TX_DATA_DEL14_reg_n_0_[37] ;
  wire \TX_DATA_DEL14_reg_n_0_[38] ;
  wire \TX_DATA_DEL14_reg_n_0_[39] ;
  wire \TX_DATA_DEL14_reg_n_0_[3] ;
  wire \TX_DATA_DEL14_reg_n_0_[40] ;
  wire \TX_DATA_DEL14_reg_n_0_[41] ;
  wire \TX_DATA_DEL14_reg_n_0_[42] ;
  wire \TX_DATA_DEL14_reg_n_0_[43] ;
  wire \TX_DATA_DEL14_reg_n_0_[44] ;
  wire \TX_DATA_DEL14_reg_n_0_[45] ;
  wire \TX_DATA_DEL14_reg_n_0_[46] ;
  wire \TX_DATA_DEL14_reg_n_0_[47] ;
  wire \TX_DATA_DEL14_reg_n_0_[48] ;
  wire \TX_DATA_DEL14_reg_n_0_[49] ;
  wire \TX_DATA_DEL14_reg_n_0_[4] ;
  wire \TX_DATA_DEL14_reg_n_0_[50] ;
  wire \TX_DATA_DEL14_reg_n_0_[51] ;
  wire \TX_DATA_DEL14_reg_n_0_[52] ;
  wire \TX_DATA_DEL14_reg_n_0_[53] ;
  wire \TX_DATA_DEL14_reg_n_0_[54] ;
  wire \TX_DATA_DEL14_reg_n_0_[55] ;
  wire \TX_DATA_DEL14_reg_n_0_[56] ;
  wire \TX_DATA_DEL14_reg_n_0_[57] ;
  wire \TX_DATA_DEL14_reg_n_0_[58] ;
  wire \TX_DATA_DEL14_reg_n_0_[59] ;
  wire \TX_DATA_DEL14_reg_n_0_[5] ;
  wire \TX_DATA_DEL14_reg_n_0_[60] ;
  wire \TX_DATA_DEL14_reg_n_0_[61] ;
  wire \TX_DATA_DEL14_reg_n_0_[62] ;
  wire \TX_DATA_DEL14_reg_n_0_[63] ;
  wire \TX_DATA_DEL14_reg_n_0_[6] ;
  wire \TX_DATA_DEL14_reg_n_0_[7] ;
  wire \TX_DATA_DEL14_reg_n_0_[8] ;
  wire \TX_DATA_DEL14_reg_n_0_[9] ;
  wire [63:0]TX_DATA_DEL15;
  wire [63:0]TX_DATA_DEL2;
  wire TX_DATA_REG0;
  wire \TX_DATA_REG[0]_i_1_n_0 ;
  wire \TX_DATA_REG[12]_i_2_n_0 ;
  wire \TX_DATA_REG[14]_i_2_n_0 ;
  wire \TX_DATA_REG[1]_i_1_n_0 ;
  wire \TX_DATA_REG[56]_i_2_n_0 ;
  wire \TX_DATA_REG[60]_i_2_n_0 ;
  wire \TX_DATA_REG[63]_i_4_n_0 ;
  wire \TX_DATA_REG[63]_i_6_n_0 ;
  wire \TX_DATA_REG[9]_i_2_n_0 ;
  wire \TX_DATA_REG_reg_n_0_[0] ;
  wire \TX_DATA_REG_reg_n_0_[10] ;
  wire \TX_DATA_REG_reg_n_0_[11] ;
  wire \TX_DATA_REG_reg_n_0_[12] ;
  wire \TX_DATA_REG_reg_n_0_[13] ;
  wire \TX_DATA_REG_reg_n_0_[14] ;
  wire \TX_DATA_REG_reg_n_0_[15] ;
  wire \TX_DATA_REG_reg_n_0_[16] ;
  wire \TX_DATA_REG_reg_n_0_[17] ;
  wire \TX_DATA_REG_reg_n_0_[18] ;
  wire \TX_DATA_REG_reg_n_0_[19] ;
  wire \TX_DATA_REG_reg_n_0_[1] ;
  wire \TX_DATA_REG_reg_n_0_[20] ;
  wire \TX_DATA_REG_reg_n_0_[21] ;
  wire \TX_DATA_REG_reg_n_0_[22] ;
  wire \TX_DATA_REG_reg_n_0_[23] ;
  wire \TX_DATA_REG_reg_n_0_[24] ;
  wire \TX_DATA_REG_reg_n_0_[25] ;
  wire \TX_DATA_REG_reg_n_0_[26] ;
  wire \TX_DATA_REG_reg_n_0_[27] ;
  wire \TX_DATA_REG_reg_n_0_[28] ;
  wire \TX_DATA_REG_reg_n_0_[29] ;
  wire \TX_DATA_REG_reg_n_0_[2] ;
  wire \TX_DATA_REG_reg_n_0_[30] ;
  wire \TX_DATA_REG_reg_n_0_[31] ;
  wire \TX_DATA_REG_reg_n_0_[32] ;
  wire \TX_DATA_REG_reg_n_0_[33] ;
  wire \TX_DATA_REG_reg_n_0_[34] ;
  wire \TX_DATA_REG_reg_n_0_[35] ;
  wire \TX_DATA_REG_reg_n_0_[36] ;
  wire \TX_DATA_REG_reg_n_0_[37] ;
  wire \TX_DATA_REG_reg_n_0_[38] ;
  wire \TX_DATA_REG_reg_n_0_[39] ;
  wire \TX_DATA_REG_reg_n_0_[3] ;
  wire \TX_DATA_REG_reg_n_0_[40] ;
  wire \TX_DATA_REG_reg_n_0_[41] ;
  wire \TX_DATA_REG_reg_n_0_[42] ;
  wire \TX_DATA_REG_reg_n_0_[43] ;
  wire \TX_DATA_REG_reg_n_0_[44] ;
  wire \TX_DATA_REG_reg_n_0_[45] ;
  wire \TX_DATA_REG_reg_n_0_[46] ;
  wire \TX_DATA_REG_reg_n_0_[47] ;
  wire \TX_DATA_REG_reg_n_0_[48] ;
  wire \TX_DATA_REG_reg_n_0_[49] ;
  wire \TX_DATA_REG_reg_n_0_[4] ;
  wire \TX_DATA_REG_reg_n_0_[50] ;
  wire \TX_DATA_REG_reg_n_0_[51] ;
  wire \TX_DATA_REG_reg_n_0_[52] ;
  wire \TX_DATA_REG_reg_n_0_[53] ;
  wire \TX_DATA_REG_reg_n_0_[54] ;
  wire \TX_DATA_REG_reg_n_0_[55] ;
  wire \TX_DATA_REG_reg_n_0_[56] ;
  wire \TX_DATA_REG_reg_n_0_[57] ;
  wire \TX_DATA_REG_reg_n_0_[58] ;
  wire \TX_DATA_REG_reg_n_0_[59] ;
  wire \TX_DATA_REG_reg_n_0_[5] ;
  wire \TX_DATA_REG_reg_n_0_[60] ;
  wire \TX_DATA_REG_reg_n_0_[61] ;
  wire \TX_DATA_REG_reg_n_0_[62] ;
  wire \TX_DATA_REG_reg_n_0_[63] ;
  wire \TX_DATA_REG_reg_n_0_[6] ;
  wire \TX_DATA_REG_reg_n_0_[7] ;
  wire \TX_DATA_REG_reg_n_0_[8] ;
  wire \TX_DATA_REG_reg_n_0_[9] ;
  wire [7:0]TX_DATA_VALID_DEL1;
  wire \TX_DATA_VALID_DEL11_reg[0]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[1]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[2]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[3]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[4]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[5]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[6]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL11_reg[7]_srl9_activity_blocks_c_7_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[0]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[1]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[2]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[3]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[4]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[5]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[6]_activity_blocks_c_8_n_0 ;
  wire \TX_DATA_VALID_DEL12_reg[7]_activity_blocks_c_8_n_0 ;
  wire [7:7]TX_DATA_VALID_DEL13;
  wire [6:0]TX_DATA_VALID_DEL13__0;
  wire [7:0]TX_DATA_VALID_DEL14;
  wire \TX_DATA_VALID_DEL14[0]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[0]_i_2_n_0 ;
  wire \TX_DATA_VALID_DEL14[1]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[1]_i_2_n_0 ;
  wire \TX_DATA_VALID_DEL14[2]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[2]_i_2_n_0 ;
  wire \TX_DATA_VALID_DEL14[3]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[4]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[5]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[5]_i_2_n_0 ;
  wire \TX_DATA_VALID_DEL14[6]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[6]_i_2_n_0 ;
  wire \TX_DATA_VALID_DEL14[6]_i_3_n_0 ;
  wire \TX_DATA_VALID_DEL14[7]_i_1_n_0 ;
  wire \TX_DATA_VALID_DEL14[7]_i_2_n_0 ;
  wire \TX_DATA_VALID_DEL14[7]_i_3_n_0 ;
  wire \TX_DATA_VALID_DEL14[7]_i_4_n_0 ;
  wire [7:0]TX_DATA_VALID_DEL15;
  wire [7:0]TX_DATA_VALID_DEL2;
  wire [63:0]TX_DATA_VALID_DELAY;
  wire [7:0]\TX_DATA_VALID_REG_reg[7]_0 ;
  wire \TX_DATA_VALID_REG_reg_n_0_[0] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[1] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[2] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[3] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[4] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[5] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[6] ;
  wire \TX_DATA_VALID_REG_reg_n_0_[7] ;
  wire TX_STATS_VALID;
  wire U_ACK_CNT_n_1;
  wire U_ACK_CNT_n_10;
  wire U_ACK_CNT_n_11;
  wire U_ACK_CNT_n_12;
  wire U_ACK_CNT_n_13;
  wire U_ACK_CNT_n_16;
  wire U_ACK_CNT_n_17;
  wire U_ACK_CNT_n_18;
  wire U_ACK_CNT_n_19;
  wire U_ACK_CNT_n_2;
  wire U_ACK_CNT_n_20;
  wire U_ACK_CNT_n_21;
  wire U_ACK_CNT_n_22;
  wire U_ACK_CNT_n_24;
  wire U_ACK_CNT_n_25;
  wire U_ACK_CNT_n_26;
  wire U_ACK_CNT_n_27;
  wire U_ACK_CNT_n_28;
  wire U_ACK_CNT_n_29;
  wire U_ACK_CNT_n_3;
  wire U_ACK_CNT_n_30;
  wire U_ACK_CNT_n_31;
  wire U_ACK_CNT_n_32;
  wire U_ACK_CNT_n_33;
  wire U_ACK_CNT_n_34;
  wire U_ACK_CNT_n_35;
  wire U_ACK_CNT_n_36;
  wire U_ACK_CNT_n_37;
  wire U_ACK_CNT_n_38;
  wire U_ACK_CNT_n_39;
  wire U_ACK_CNT_n_4;
  wire U_ACK_CNT_n_5;
  wire U_ACK_CNT_n_6;
  wire U_ACK_CNT_n_7;
  wire U_ACK_CNT_n_8;
  wire U_ACK_CNT_n_9;
  wire U_CRC8_n_0;
  wire U_CRC8_n_1;
  wire U_CRC8_n_10;
  wire U_CRC8_n_11;
  wire U_CRC8_n_12;
  wire U_CRC8_n_13;
  wire U_CRC8_n_14;
  wire U_CRC8_n_15;
  wire U_CRC8_n_16;
  wire U_CRC8_n_17;
  wire U_CRC8_n_18;
  wire U_CRC8_n_19;
  wire U_CRC8_n_2;
  wire U_CRC8_n_20;
  wire U_CRC8_n_21;
  wire U_CRC8_n_22;
  wire U_CRC8_n_23;
  wire U_CRC8_n_24;
  wire U_CRC8_n_25;
  wire U_CRC8_n_26;
  wire U_CRC8_n_27;
  wire U_CRC8_n_28;
  wire U_CRC8_n_29;
  wire U_CRC8_n_3;
  wire U_CRC8_n_30;
  wire U_CRC8_n_31;
  wire U_CRC8_n_32;
  wire U_CRC8_n_33;
  wire U_CRC8_n_34;
  wire U_CRC8_n_35;
  wire U_CRC8_n_36;
  wire U_CRC8_n_37;
  wire U_CRC8_n_38;
  wire U_CRC8_n_39;
  wire U_CRC8_n_4;
  wire U_CRC8_n_40;
  wire U_CRC8_n_41;
  wire U_CRC8_n_42;
  wire U_CRC8_n_43;
  wire U_CRC8_n_44;
  wire U_CRC8_n_45;
  wire U_CRC8_n_46;
  wire U_CRC8_n_47;
  wire U_CRC8_n_48;
  wire U_CRC8_n_49;
  wire U_CRC8_n_5;
  wire U_CRC8_n_50;
  wire U_CRC8_n_51;
  wire U_CRC8_n_52;
  wire U_CRC8_n_53;
  wire U_CRC8_n_54;
  wire U_CRC8_n_55;
  wire U_CRC8_n_56;
  wire U_CRC8_n_57;
  wire U_CRC8_n_58;
  wire U_CRC8_n_59;
  wire U_CRC8_n_6;
  wire U_CRC8_n_60;
  wire U_CRC8_n_61;
  wire U_CRC8_n_62;
  wire U_CRC8_n_63;
  wire U_CRC8_n_64;
  wire U_CRC8_n_65;
  wire U_CRC8_n_66;
  wire U_CRC8_n_67;
  wire U_CRC8_n_68;
  wire U_CRC8_n_69;
  wire U_CRC8_n_7;
  wire U_CRC8_n_70;
  wire U_CRC8_n_71;
  wire U_CRC8_n_72;
  wire U_CRC8_n_73;
  wire U_CRC8_n_74;
  wire U_CRC8_n_75;
  wire U_CRC8_n_76;
  wire U_CRC8_n_77;
  wire U_CRC8_n_78;
  wire U_CRC8_n_79;
  wire U_CRC8_n_8;
  wire U_CRC8_n_80;
  wire U_CRC8_n_81;
  wire U_CRC8_n_82;
  wire U_CRC8_n_83;
  wire U_CRC8_n_84;
  wire U_CRC8_n_85;
  wire U_CRC8_n_86;
  wire U_CRC8_n_87;
  wire U_CRC8_n_88;
  wire U_CRC8_n_9;
  wire U_byte_count_module_n_100;
  wire U_byte_count_module_n_101;
  wire U_byte_count_module_n_102;
  wire U_byte_count_module_n_103;
  wire U_byte_count_module_n_104;
  wire U_byte_count_module_n_105;
  wire U_byte_count_module_n_107;
  wire U_byte_count_module_n_28;
  wire U_byte_count_module_n_29;
  wire U_byte_count_module_n_30;
  wire U_byte_count_module_n_31;
  wire U_byte_count_module_n_32;
  wire U_byte_count_module_n_33;
  wire U_byte_count_module_n_34;
  wire U_byte_count_module_n_35;
  wire U_byte_count_module_n_36;
  wire U_byte_count_module_n_37;
  wire U_byte_count_module_n_38;
  wire U_byte_count_module_n_39;
  wire U_byte_count_module_n_40;
  wire U_byte_count_module_n_41;
  wire U_byte_count_module_n_42;
  wire U_byte_count_module_n_43;
  wire U_byte_count_module_n_45;
  wire U_byte_count_module_n_46;
  wire U_byte_count_module_n_47;
  wire U_byte_count_module_n_48;
  wire U_byte_count_module_n_49;
  wire U_byte_count_module_n_50;
  wire U_byte_count_module_n_51;
  wire U_byte_count_module_n_52;
  wire U_byte_count_module_n_53;
  wire U_byte_count_module_n_54;
  wire U_byte_count_module_n_55;
  wire U_byte_count_module_n_56;
  wire U_byte_count_module_n_57;
  wire U_byte_count_module_n_58;
  wire U_byte_count_module_n_59;
  wire U_byte_count_module_n_60;
  wire U_byte_count_module_n_61;
  wire U_byte_count_module_n_62;
  wire U_byte_count_module_n_63;
  wire U_byte_count_module_n_64;
  wire U_byte_count_module_n_65;
  wire U_byte_count_module_n_66;
  wire U_byte_count_module_n_67;
  wire U_byte_count_module_n_68;
  wire U_byte_count_module_n_69;
  wire U_byte_count_module_n_70;
  wire U_byte_count_module_n_71;
  wire U_byte_count_module_n_72;
  wire U_byte_count_module_n_73;
  wire U_byte_count_module_n_74;
  wire U_byte_count_module_n_75;
  wire U_byte_count_module_n_76;
  wire U_byte_count_module_n_77;
  wire U_byte_count_module_n_78;
  wire U_byte_count_module_n_79;
  wire U_byte_count_module_n_80;
  wire U_byte_count_module_n_81;
  wire U_byte_count_module_n_82;
  wire U_byte_count_module_n_83;
  wire U_byte_count_module_n_84;
  wire U_byte_count_module_n_85;
  wire U_byte_count_module_n_86;
  wire U_byte_count_module_n_87;
  wire U_byte_count_module_n_88;
  wire U_byte_count_module_n_89;
  wire U_byte_count_module_n_90;
  wire U_byte_count_module_n_91;
  wire U_byte_count_module_n_92;
  wire U_byte_count_module_n_93;
  wire U_byte_count_module_n_94;
  wire U_byte_count_module_n_95;
  wire U_byte_count_module_n_96;
  wire U_byte_count_module_n_97;
  wire U_byte_count_module_n_98;
  wire U_byte_count_module_n_99;
  wire activity_blocks_gate__0_n_0;
  wire activity_blocks_gate__10_n_0;
  wire activity_blocks_gate__11_n_0;
  wire activity_blocks_gate__12_n_0;
  wire activity_blocks_gate__13_n_0;
  wire activity_blocks_gate__14_n_0;
  wire activity_blocks_gate__15_n_0;
  wire activity_blocks_gate__16_n_0;
  wire activity_blocks_gate__17_n_0;
  wire activity_blocks_gate__18_n_0;
  wire activity_blocks_gate__19_n_0;
  wire activity_blocks_gate__1_n_0;
  wire activity_blocks_gate__20_n_0;
  wire activity_blocks_gate__21_n_0;
  wire activity_blocks_gate__22_n_0;
  wire activity_blocks_gate__23_n_0;
  wire activity_blocks_gate__24_n_0;
  wire activity_blocks_gate__25_n_0;
  wire activity_blocks_gate__26_n_0;
  wire activity_blocks_gate__27_n_0;
  wire activity_blocks_gate__28_n_0;
  wire activity_blocks_gate__29_n_0;
  wire activity_blocks_gate__2_n_0;
  wire activity_blocks_gate__30_n_0;
  wire activity_blocks_gate__31_n_0;
  wire activity_blocks_gate__32_n_0;
  wire activity_blocks_gate__33_n_0;
  wire activity_blocks_gate__34_n_0;
  wire activity_blocks_gate__35_n_0;
  wire activity_blocks_gate__36_n_0;
  wire activity_blocks_gate__37_n_0;
  wire activity_blocks_gate__38_n_0;
  wire activity_blocks_gate__39_n_0;
  wire activity_blocks_gate__3_n_0;
  wire activity_blocks_gate__40_n_0;
  wire activity_blocks_gate__41_n_0;
  wire activity_blocks_gate__42_n_0;
  wire activity_blocks_gate__43_n_0;
  wire activity_blocks_gate__44_n_0;
  wire activity_blocks_gate__45_n_0;
  wire activity_blocks_gate__46_n_0;
  wire activity_blocks_gate__47_n_0;
  wire activity_blocks_gate__48_n_0;
  wire activity_blocks_gate__49_n_0;
  wire activity_blocks_gate__4_n_0;
  wire activity_blocks_gate__50_n_0;
  wire activity_blocks_gate__51_n_0;
  wire activity_blocks_gate__52_n_0;
  wire activity_blocks_gate__53_n_0;
  wire activity_blocks_gate__54_n_0;
  wire activity_blocks_gate__55_n_0;
  wire activity_blocks_gate__56_n_0;
  wire activity_blocks_gate__57_n_0;
  wire activity_blocks_gate__58_n_0;
  wire activity_blocks_gate__59_n_0;
  wire activity_blocks_gate__5_n_0;
  wire activity_blocks_gate__60_n_0;
  wire activity_blocks_gate__61_n_0;
  wire activity_blocks_gate__62_n_0;
  wire activity_blocks_gate__63_n_0;
  wire activity_blocks_gate__64_n_0;
  wire activity_blocks_gate__65_n_0;
  wire activity_blocks_gate__66_n_0;
  wire activity_blocks_gate__67_n_0;
  wire activity_blocks_gate__68_n_0;
  wire activity_blocks_gate__69_n_0;
  wire activity_blocks_gate__6_n_0;
  wire activity_blocks_gate__70_n_0;
  wire activity_blocks_gate__71_n_0;
  wire activity_blocks_gate__7_n_0;
  wire activity_blocks_gate__8_n_0;
  wire activity_blocks_gate__9_n_0;
  wire activity_blocks_gate_n_0;
  wire append_end_frame;
  wire \append_reg_reg[8]_srl9_activity_blocks_c_7_n_0 ;
  wire \append_reg_reg[9]_activity_blocks_c_8_n_0 ;
  wire append_start_pause;
  wire append_start_pause0;
  wire apply_pause_delay;
  wire apply_pause_delay_reg_0;
  wire apply_pause_delay_reg_n_0;
  wire [15:2]byte_count_reg;
  wire \byte_count_stat_reg_n_0_[0] ;
  wire \byte_count_stat_reg_n_0_[10] ;
  wire \byte_count_stat_reg_n_0_[11] ;
  wire \byte_count_stat_reg_n_0_[12] ;
  wire \byte_count_stat_reg_n_0_[13] ;
  wire \byte_count_stat_reg_n_0_[1] ;
  wire \byte_count_stat_reg_n_0_[2] ;
  wire \byte_count_stat_reg_n_0_[3] ;
  wire \byte_count_stat_reg_n_0_[4] ;
  wire \byte_count_stat_reg_n_0_[5] ;
  wire \byte_count_stat_reg_n_0_[6] ;
  wire \byte_count_stat_reg_n_0_[7] ;
  wire \byte_count_stat_reg_n_0_[8] ;
  wire \byte_count_stat_reg_n_0_[9] ;
  wire clk_i;
  wire fcs_enabled_int;
  wire \final_byte_count[10]_i_2_n_0 ;
  wire \final_byte_count[12]_i_2_n_0 ;
  wire \final_byte_count[13]_i_2_n_0 ;
  wire \final_byte_count[13]_i_3_n_0 ;
  wire \final_byte_count[15]_i_3_n_0 ;
  wire \final_byte_count[3]_i_2_n_0 ;
  wire \final_byte_count[4]_i_2_n_0 ;
  wire \final_byte_count[5]_i_3_n_0 ;
  wire \final_byte_count[7]_i_2_n_0 ;
  wire \final_byte_count[8]_i_2_n_0 ;
  wire \final_byte_count[9]_i_2_n_0 ;
  wire [13:0]final_byte_count_reg;
  wire [15:14]final_byte_count_reg__0;
  wire frame_start_del;
  wire insert_error1__0;
  wire insert_error_i_10_n_0;
  wire insert_error_i_11_n_0;
  wire insert_error_i_12_n_0;
  wire insert_error_i_13_n_0;
  wire insert_error_i_14_n_0;
  wire insert_error_i_15_n_0;
  wire insert_error_i_16_n_0;
  wire insert_error_i_17_n_0;
  wire insert_error_i_18_n_0;
  wire insert_error_i_19_n_0;
  wire insert_error_i_1_n_0;
  wire insert_error_i_20_n_0;
  wire insert_error_i_21_n_0;
  wire insert_error_i_22_n_0;
  wire insert_error_i_23_n_0;
  wire insert_error_i_24_n_0;
  wire insert_error_i_25_n_0;
  wire insert_error_i_26_n_0;
  wire insert_error_i_27_n_0;
  wire insert_error_i_28_n_0;
  wire insert_error_i_29_n_0;
  wire insert_error_i_2_n_0;
  wire insert_error_i_30_n_0;
  wire insert_error_i_31_n_0;
  wire insert_error_i_3_n_0;
  wire insert_error_i_4_n_0;
  wire insert_error_i_5_n_0;
  wire insert_error_i_6_n_0;
  wire insert_error_i_8_n_0;
  wire insert_error_i_9_n_0;
  wire insert_error_reg_i_7_n_1;
  wire insert_error_reg_i_7_n_2;
  wire insert_error_reg_i_7_n_3;
  wire insert_error_reg_i_7_n_4;
  wire insert_error_reg_i_7_n_5;
  wire insert_error_reg_i_7_n_6;
  wire insert_error_reg_i_7_n_7;
  wire [15:0]length_register;
  wire length_register0;
  wire load_CRC8;
  wire load_CRC80;
  wire load_final_CRC_reg_0;
  wire out;
  wire [3:1]p_0_in__0;
  wire [15:0]p_0_in__2;
  wire pause_frame_counter0;
  wire \pause_frame_counter[0]_i_1_n_0 ;
  wire [3:0]pause_frame_counter_reg;
  wire read_ifg_int;
  wire reset_err_pause;
  wire reset_err_pause0;
  wire reset_tx_int;
  wire rst_i;
  wire set_pause_stats;
  wire set_pause_stats_i_1_n_0;
  wire [60:0]shift_pause_data;
  wire \shift_pause_data[0]_i_1_n_0 ;
  wire \shift_pause_data[10]_i_1_n_0 ;
  wire \shift_pause_data[11]_i_1_n_0 ;
  wire \shift_pause_data[12]_i_1_n_0 ;
  wire \shift_pause_data[13]_i_1_n_0 ;
  wire \shift_pause_data[14]_i_1_n_0 ;
  wire \shift_pause_data[15]_i_1_n_0 ;
  wire \shift_pause_data[1]_i_1_n_0 ;
  wire \shift_pause_data[2]_i_1_n_0 ;
  wire \shift_pause_data[3]_i_1_n_0 ;
  wire \shift_pause_data[4]_i_1_n_0 ;
  wire \shift_pause_data[56]_i_1_n_0 ;
  wire \shift_pause_data[56]_i_2_n_0 ;
  wire \shift_pause_data[5]_i_1_n_0 ;
  wire \shift_pause_data[60]_i_1_n_0 ;
  wire \shift_pause_data[6]_i_1_n_0 ;
  wire \shift_pause_data[7]_i_1_n_0 ;
  wire \shift_pause_data[8]_i_1_n_0 ;
  wire \shift_pause_data[9]_i_1_n_0 ;
  wire [4:0]shift_pause_valid;
  wire \shift_pause_valid[0]_i_1_n_0 ;
  wire \shift_pause_valid[4]_i_1_n_0 ;
  wire [4:0]shift_pause_valid_del;
  wire start_CRC8;
  wire [15:0]store_pause_frame;
  wire \store_tx_data[0]_i_1_n_0 ;
  wire \store_tx_data[10]_i_1_n_0 ;
  wire \store_tx_data[11]_i_1_n_0 ;
  wire \store_tx_data[12]_i_1_n_0 ;
  wire \store_tx_data[13]_i_1_n_0 ;
  wire \store_tx_data[14]_i_1_n_0 ;
  wire \store_tx_data[15]_i_1_n_0 ;
  wire \store_tx_data[16]_i_1_n_0 ;
  wire \store_tx_data[17]_i_1_n_0 ;
  wire \store_tx_data[18]_i_1_n_0 ;
  wire \store_tx_data[19]_i_1_n_0 ;
  wire \store_tx_data[1]_i_1_n_0 ;
  wire \store_tx_data[20]_i_1_n_0 ;
  wire \store_tx_data[21]_i_1_n_0 ;
  wire \store_tx_data[22]_i_1_n_0 ;
  wire \store_tx_data[23]_i_1_n_0 ;
  wire \store_tx_data[24]_i_1_n_0 ;
  wire \store_tx_data[25]_i_1_n_0 ;
  wire \store_tx_data[26]_i_1_n_0 ;
  wire \store_tx_data[27]_i_1_n_0 ;
  wire \store_tx_data[28]_i_1_n_0 ;
  wire \store_tx_data[29]_i_1_n_0 ;
  wire \store_tx_data[2]_i_1_n_0 ;
  wire \store_tx_data[30]_i_1_n_0 ;
  wire \store_tx_data[31]_i_1_n_0 ;
  wire \store_tx_data[32]_i_1_n_0 ;
  wire \store_tx_data[33]_i_1_n_0 ;
  wire \store_tx_data[34]_i_1_n_0 ;
  wire \store_tx_data[35]_i_1_n_0 ;
  wire \store_tx_data[36]_i_1_n_0 ;
  wire \store_tx_data[37]_i_1_n_0 ;
  wire \store_tx_data[38]_i_1_n_0 ;
  wire \store_tx_data[39]_i_1_n_0 ;
  wire \store_tx_data[3]_i_1_n_0 ;
  wire \store_tx_data[40]_i_1_n_0 ;
  wire \store_tx_data[41]_i_1_n_0 ;
  wire \store_tx_data[42]_i_1_n_0 ;
  wire \store_tx_data[43]_i_1_n_0 ;
  wire \store_tx_data[44]_i_1_n_0 ;
  wire \store_tx_data[45]_i_1_n_0 ;
  wire \store_tx_data[46]_i_1_n_0 ;
  wire \store_tx_data[47]_i_1_n_0 ;
  wire \store_tx_data[48]_i_1_n_0 ;
  wire \store_tx_data[49]_i_1_n_0 ;
  wire \store_tx_data[4]_i_1_n_0 ;
  wire \store_tx_data[50]_i_1_n_0 ;
  wire \store_tx_data[51]_i_1_n_0 ;
  wire \store_tx_data[52]_i_1_n_0 ;
  wire \store_tx_data[53]_i_1_n_0 ;
  wire \store_tx_data[54]_i_1_n_0 ;
  wire \store_tx_data[55]_i_1_n_0 ;
  wire \store_tx_data[5]_i_1_n_0 ;
  wire \store_tx_data[6]_i_1_n_0 ;
  wire \store_tx_data[7]_i_1_n_0 ;
  wire \store_tx_data[8]_i_1_n_0 ;
  wire \store_tx_data[9]_i_1_n_0 ;
  wire \store_tx_data_reg_n_0_[0] ;
  wire \store_tx_data_reg_n_0_[10] ;
  wire \store_tx_data_reg_n_0_[11] ;
  wire \store_tx_data_reg_n_0_[12] ;
  wire \store_tx_data_reg_n_0_[13] ;
  wire \store_tx_data_reg_n_0_[14] ;
  wire \store_tx_data_reg_n_0_[15] ;
  wire \store_tx_data_reg_n_0_[16] ;
  wire \store_tx_data_reg_n_0_[17] ;
  wire \store_tx_data_reg_n_0_[18] ;
  wire \store_tx_data_reg_n_0_[19] ;
  wire \store_tx_data_reg_n_0_[1] ;
  wire \store_tx_data_reg_n_0_[20] ;
  wire \store_tx_data_reg_n_0_[21] ;
  wire \store_tx_data_reg_n_0_[22] ;
  wire \store_tx_data_reg_n_0_[23] ;
  wire \store_tx_data_reg_n_0_[24] ;
  wire \store_tx_data_reg_n_0_[25] ;
  wire \store_tx_data_reg_n_0_[26] ;
  wire \store_tx_data_reg_n_0_[27] ;
  wire \store_tx_data_reg_n_0_[28] ;
  wire \store_tx_data_reg_n_0_[29] ;
  wire \store_tx_data_reg_n_0_[2] ;
  wire \store_tx_data_reg_n_0_[30] ;
  wire \store_tx_data_reg_n_0_[31] ;
  wire \store_tx_data_reg_n_0_[32] ;
  wire \store_tx_data_reg_n_0_[33] ;
  wire \store_tx_data_reg_n_0_[34] ;
  wire \store_tx_data_reg_n_0_[35] ;
  wire \store_tx_data_reg_n_0_[36] ;
  wire \store_tx_data_reg_n_0_[37] ;
  wire \store_tx_data_reg_n_0_[38] ;
  wire \store_tx_data_reg_n_0_[39] ;
  wire \store_tx_data_reg_n_0_[3] ;
  wire \store_tx_data_reg_n_0_[40] ;
  wire \store_tx_data_reg_n_0_[41] ;
  wire \store_tx_data_reg_n_0_[42] ;
  wire \store_tx_data_reg_n_0_[43] ;
  wire \store_tx_data_reg_n_0_[44] ;
  wire \store_tx_data_reg_n_0_[45] ;
  wire \store_tx_data_reg_n_0_[46] ;
  wire \store_tx_data_reg_n_0_[47] ;
  wire \store_tx_data_reg_n_0_[48] ;
  wire \store_tx_data_reg_n_0_[49] ;
  wire \store_tx_data_reg_n_0_[4] ;
  wire \store_tx_data_reg_n_0_[50] ;
  wire \store_tx_data_reg_n_0_[51] ;
  wire \store_tx_data_reg_n_0_[52] ;
  wire \store_tx_data_reg_n_0_[53] ;
  wire \store_tx_data_reg_n_0_[54] ;
  wire \store_tx_data_reg_n_0_[55] ;
  wire \store_tx_data_reg_n_0_[56] ;
  wire \store_tx_data_reg_n_0_[57] ;
  wire \store_tx_data_reg_n_0_[58] ;
  wire \store_tx_data_reg_n_0_[59] ;
  wire \store_tx_data_reg_n_0_[5] ;
  wire \store_tx_data_reg_n_0_[60] ;
  wire \store_tx_data_reg_n_0_[61] ;
  wire \store_tx_data_reg_n_0_[62] ;
  wire \store_tx_data_reg_n_0_[63] ;
  wire \store_tx_data_reg_n_0_[6] ;
  wire \store_tx_data_reg_n_0_[7] ;
  wire \store_tx_data_reg_n_0_[8] ;
  wire \store_tx_data_reg_n_0_[9] ;
  wire \store_tx_data_valid[0]_i_1_n_0 ;
  wire \store_tx_data_valid[1]_i_1_n_0 ;
  wire \store_tx_data_valid[2]_i_1_n_0 ;
  wire \store_tx_data_valid[3]_i_1_n_0 ;
  wire \store_tx_data_valid[4]_i_1_n_0 ;
  wire \store_tx_data_valid[5]_i_1_n_0 ;
  wire \store_tx_data_valid[6]_i_1_n_0 ;
  wire \store_tx_data_valid_reg_n_0_[0] ;
  wire \store_tx_data_valid_reg_n_0_[1] ;
  wire \store_tx_data_valid_reg_n_0_[2] ;
  wire \store_tx_data_valid_reg_n_0_[3] ;
  wire \store_tx_data_valid_reg_n_0_[4] ;
  wire \store_tx_data_valid_reg_n_0_[5] ;
  wire \store_tx_data_valid_reg_n_0_[6] ;
  wire \store_tx_data_valid_reg_n_0_[7] ;
  wire transmit_pause_frame_del;
  wire transmit_pause_frame_del2;
  wire transmit_pause_frame_del3;
  wire transmit_pause_frame_i_1_n_0;
  wire transmit_pause_frame_reg_n_0;
  wire transmit_pause_frame_valid;
  wire transmit_pause_frame_valid0;
  wire [7:0]tx_data_int;
  wire \tx_data_int[7]_i_1_n_0 ;
  wire tx_undderrun_int;
  wire tx_undderrun_int_i_1_n_0;
  wire tx_undderrun_int_reg_0;
  wire [3:3]txstatplus_int;
  wire [18:1]txstatplus_int0_out;
  wire \txstatplus_int[18]_i_1_n_0 ;
  wire \txstatplus_int[19]_i_1_n_0 ;
  wire \txstatplus_int[24]_i_1_n_0 ;
  wire \txstatplus_int[3]_i_1_n_0 ;
  wire \txstatplus_int_reg_n_0_[10] ;
  wire \txstatplus_int_reg_n_0_[11] ;
  wire \txstatplus_int_reg_n_0_[12] ;
  wire \txstatplus_int_reg_n_0_[13] ;
  wire \txstatplus_int_reg_n_0_[14] ;
  wire \txstatplus_int_reg_n_0_[15] ;
  wire \txstatplus_int_reg_n_0_[16] ;
  wire \txstatplus_int_reg_n_0_[17] ;
  wire \txstatplus_int_reg_n_0_[18] ;
  wire \txstatplus_int_reg_n_0_[19] ;
  wire \txstatplus_int_reg_n_0_[1] ;
  wire \txstatplus_int_reg_n_0_[24] ;
  wire \txstatplus_int_reg_n_0_[2] ;
  wire \txstatplus_int_reg_n_0_[3] ;
  wire \txstatplus_int_reg_n_0_[4] ;
  wire \txstatplus_int_reg_n_0_[5] ;
  wire \txstatplus_int_reg_n_0_[6] ;
  wire \txstatplus_int_reg_n_0_[7] ;
  wire \txstatplus_int_reg_n_0_[8] ;
  wire \txstatplus_int_reg_n_0_[9] ;
  wire vlan_enabled_int;
  wire [7:0]NLW_insert_error_reg_i_7_O_UNCONNECTED;

  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[0]_i_1 
       (.I0(store_pause_frame[0]),
        .I1(\DELAY_ACK_reg[7]_0 [0]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair450" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[10]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[10]),
        .O(\DELAY_ACK[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair451" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[11]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[11]),
        .O(\DELAY_ACK[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair452" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[12]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[12]),
        .O(\DELAY_ACK[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair453" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[13]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[13]),
        .O(\DELAY_ACK[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair470" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[14]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[14]),
        .O(\DELAY_ACK[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \DELAY_ACK[15]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(read_ifg_int),
        .O(\DELAY_ACK[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[15]_i_2 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[15]),
        .O(\DELAY_ACK[15]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair453" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[1]_i_1 
       (.I0(store_pause_frame[1]),
        .I1(\DELAY_ACK_reg[7]_0 [1]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair452" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[2]_i_1 
       (.I0(store_pause_frame[2]),
        .I1(\DELAY_ACK_reg[7]_0 [2]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair451" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[3]_i_1 
       (.I0(store_pause_frame[3]),
        .I1(\DELAY_ACK_reg[7]_0 [3]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair450" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[4]_i_1 
       (.I0(store_pause_frame[4]),
        .I1(\DELAY_ACK_reg[7]_0 [4]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair449" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[5]_i_1 
       (.I0(store_pause_frame[5]),
        .I1(\DELAY_ACK_reg[7]_0 [5]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair470" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[6]_i_1 
       (.I0(store_pause_frame[6]),
        .I1(\DELAY_ACK_reg[7]_0 [6]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair448" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \DELAY_ACK[7]_i_1 
       (.I0(store_pause_frame[7]),
        .I1(\DELAY_ACK_reg[7]_0 [7]),
        .I2(apply_pause_delay_reg_n_0),
        .O(\DELAY_ACK[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair448" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[8]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[8]),
        .O(\DELAY_ACK[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair449" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \DELAY_ACK[9]_i_1 
       (.I0(apply_pause_delay_reg_n_0),
        .I1(store_pause_frame[9]),
        .O(\DELAY_ACK[9]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \DELAY_ACK_reg[0] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .D(\DELAY_ACK[0]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(DELAY_ACK[0]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[10] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[10]_i_1_n_0 ),
        .Q(DELAY_ACK[10]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[11] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[11]_i_1_n_0 ),
        .Q(DELAY_ACK[11]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[12] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[12]_i_1_n_0 ),
        .Q(DELAY_ACK[12]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[13] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[13]_i_1_n_0 ),
        .Q(DELAY_ACK[13]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[14] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[14]_i_1_n_0 ),
        .Q(DELAY_ACK[14]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[15] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[15]_i_2_n_0 ),
        .Q(DELAY_ACK[15]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[1] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[1]_i_1_n_0 ),
        .Q(DELAY_ACK[1]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[2] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[2]_i_1_n_0 ),
        .Q(DELAY_ACK[2]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[3] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[3]_i_1_n_0 ),
        .Q(DELAY_ACK[3]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[4] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[4]_i_1_n_0 ),
        .Q(DELAY_ACK[4]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[5] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[5]_i_1_n_0 ),
        .Q(DELAY_ACK[5]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[6] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[6]_i_1_n_0 ),
        .Q(DELAY_ACK[6]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[7] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[7]_i_1_n_0 ),
        .Q(DELAY_ACK[7]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[8] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[8]_i_1_n_0 ),
        .Q(DELAY_ACK[8]));
  FDCE #(
    .INIT(1'b0)) 
    \DELAY_ACK_reg[9] 
       (.C(clk_i),
        .CE(\DELAY_ACK[15]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\DELAY_ACK[9]_i_1_n_0 ),
        .Q(DELAY_ACK[9]));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    FRAME_START_i_3
       (.I0(\TX_DATA_VALID_REG_reg_n_0_[7] ),
        .I1(\TX_DATA_VALID_REG_reg_n_0_[6] ),
        .I2(\TX_DATA_VALID_REG_reg_n_0_[4] ),
        .I3(\TX_DATA_VALID_REG_reg_n_0_[5] ),
        .I4(FRAME_START_i_4_n_0),
        .O(FRAME_START_i_3_n_0));
  (* SOFT_HLUTNM = "soft_lutpair429" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    FRAME_START_i_4
       (.I0(\TX_DATA_VALID_REG_reg_n_0_[1] ),
        .I1(\TX_DATA_VALID_REG_reg_n_0_[0] ),
        .I2(\TX_DATA_VALID_REG_reg_n_0_[3] ),
        .I3(\TX_DATA_VALID_REG_reg_n_0_[2] ),
        .O(FRAME_START_i_4_n_0));
  FDCE #(
    .INIT(1'b0)) 
    FRAME_START_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_107),
        .Q(FRAME_START));
  LUT2 #(
    .INIT(4'h6)) 
    \MAX_FRAME_SIZE[2]_i_1 
       (.I0(fcs_enabled_int),
        .I1(vlan_enabled_int),
        .O(\MAX_FRAME_SIZE[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair444" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \MAX_FRAME_SIZE[3]_i_1 
       (.I0(vlan_enabled_int),
        .I1(fcs_enabled_int),
        .O(\MAX_FRAME_SIZE[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair446" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \MAX_FRAME_SIZE[4]_i_1 
       (.I0(fcs_enabled_int),
        .I1(vlan_enabled_int),
        .O(\MAX_FRAME_SIZE[4]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \MAX_FRAME_SIZE_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\MAX_FRAME_SIZE[2]_i_1_n_0 ),
        .Q(MAX_FRAME_SIZE[2]));
  FDPE #(
    .INIT(1'b1)) 
    \MAX_FRAME_SIZE_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\MAX_FRAME_SIZE[3]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(MAX_FRAME_SIZE[3]));
  FDCE #(
    .INIT(1'b0)) 
    \MAX_FRAME_SIZE_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\MAX_FRAME_SIZE[4]_i_1_n_0 ),
        .Q(MAX_FRAME_SIZE[4]));
  (* SOFT_HLUTNM = "soft_lutpair421" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \OVERFLOW_DATA[17]_i_2 
       (.I0(TX_DATA_VALID_DEL13__0[2]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .O(\OVERFLOW_DATA[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00D5D5D500000000)) 
    \OVERFLOW_DATA[23]_i_2 
       (.I0(\OVERFLOW_DATA[31]_i_2_n_0 ),
        .I1(txstatplus_int),
        .I2(fcs_enabled_int),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[6]),
        .I5(TX_DATA_VALID_DEL13__0[4]),
        .O(\OVERFLOW_DATA[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF3AFAFAFFFFFFFFF)) 
    \OVERFLOW_DATA[25]_i_1 
       (.I0(\OVERFLOW_DATA[31]_i_2_n_0 ),
        .I1(fcs_enabled_int),
        .I2(txstatplus_int),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[6]),
        .I5(TX_DATA_VALID_DEL13__0[4]),
        .O(\OVERFLOW_DATA[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h80008CCC80008000)) 
    \OVERFLOW_DATA[31]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[4]),
        .I2(TX_DATA_VALID_DEL13__0[6]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(\OVERFLOW_DATA[31]_i_2_n_0 ),
        .I5(txstatplus_int),
        .O(\OVERFLOW_DATA[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8AFF000000000000)) 
    \OVERFLOW_DATA[31]_i_2 
       (.I0(TX_DATA_VALID_DEL13__0[4]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(TX_DATA_VALID_DEL13__0[1]),
        .I5(TX_DATA_VALID_DEL13__0[2]),
        .O(\OVERFLOW_DATA[31]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair421" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \OVERFLOW_DATA[33]_i_1 
       (.I0(fcs_enabled_int),
        .I1(txstatplus_int),
        .I2(TX_DATA_VALID_DEL13__0[2]),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .O(\OVERFLOW_DATA[33]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hAA8A)) 
    \OVERFLOW_DATA[39]_i_1 
       (.I0(\OVERFLOW_VALID[2]_i_1_n_0 ),
        .I1(fcs_enabled_int),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .O(\OVERFLOW_DATA[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair424" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \OVERFLOW_DATA[39]_i_2 
       (.I0(TX_DATA_VALID_DEL13__0[4]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[2]),
        .I3(txstatplus_int),
        .I4(fcs_enabled_int),
        .O(\OVERFLOW_DATA[39]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair424" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \OVERFLOW_DATA[8]_i_2 
       (.I0(fcs_enabled_int),
        .I1(txstatplus_int),
        .O(\OVERFLOW_DATA[8]_i_2_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[0] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_23),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[0] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[10] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_13),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[11] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_12),
        .Q(\OVERFLOW_DATA_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[12] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_11),
        .Q(\OVERFLOW_DATA_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[13] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_10),
        .Q(\OVERFLOW_DATA_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[14] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_9),
        .Q(\OVERFLOW_DATA_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[15] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_8),
        .Q(\OVERFLOW_DATA_reg_n_0_[15] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[16] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_7),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[16] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[17] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_6),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[17] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[18] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_5),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[19] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_4),
        .Q(\OVERFLOW_DATA_reg_n_0_[19] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[1] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_22),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[20] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_3),
        .Q(\OVERFLOW_DATA_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[21] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_2),
        .Q(\OVERFLOW_DATA_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[22] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_1),
        .Q(\OVERFLOW_DATA_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[23] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_0),
        .Q(\OVERFLOW_DATA_reg_n_0_[23] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[25] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(\OVERFLOW_DATA[25]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[25] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[2] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_21),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[31] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\OVERFLOW_DATA[31]_i_1_n_0 ),
        .Q(\OVERFLOW_DATA_reg_n_0_[31] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[33] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(\OVERFLOW_DATA[33]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[39] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\OVERFLOW_DATA[39]_i_2_n_0 ),
        .Q(\OVERFLOW_DATA_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[3] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_20),
        .Q(\OVERFLOW_DATA_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[4] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_19),
        .Q(\OVERFLOW_DATA_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[5] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_18),
        .Q(\OVERFLOW_DATA_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[6] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_17),
        .Q(\OVERFLOW_DATA_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_DATA_reg[7] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .CLR(rst_i),
        .D(U_CRC8_n_16),
        .Q(\OVERFLOW_DATA_reg_n_0_[7] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[8] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_15),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[8] ));
  FDPE #(
    .INIT(1'b1)) 
    \OVERFLOW_DATA_reg[9] 
       (.C(clk_i),
        .CE(\OVERFLOW_DATA[39]_i_1_n_0 ),
        .D(U_CRC8_n_14),
        .PRE(rst_i),
        .Q(\OVERFLOW_DATA_reg_n_0_[9] ));
  LUT2 #(
    .INIT(4'h8)) 
    \OVERFLOW_VALID[0]_i_1 
       (.I0(TX_DATA_VALID_DEL13__0[4]),
        .I1(fcs_enabled_int),
        .O(\OVERFLOW_VALID[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair516" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \OVERFLOW_VALID[1]_i_1 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[5]),
        .O(\OVERFLOW_VALID[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000808000C5)) 
    \OVERFLOW_VALID[2]_i_1 
       (.I0(TX_DATA_VALID_DEL13__0[2]),
        .I1(TX_DATA_VALID_DEL13__0[0]),
        .I2(TX_DATA_VALID_DEL13__0[1]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[3]),
        .I5(\OVERFLOW_VALID[2]_i_3_n_0 ),
        .O(\OVERFLOW_VALID[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair516" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \OVERFLOW_VALID[2]_i_2 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .O(\OVERFLOW_VALID[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair420" *) 
  LUT5 #(
    .INIT(32'hBBFBFFFB)) 
    \OVERFLOW_VALID[2]_i_3 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(txstatplus_int0_out[1]),
        .I2(TX_DATA_VALID_DEL13__0[6]),
        .I3(TX_DATA_VALID_DEL13__0[5]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .O(\OVERFLOW_VALID[2]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_VALID_reg[0] 
       (.C(clk_i),
        .CE(\OVERFLOW_VALID[2]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\OVERFLOW_VALID[0]_i_1_n_0 ),
        .Q(OVERFLOW_VALID__0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_VALID_reg[1] 
       (.C(clk_i),
        .CE(\OVERFLOW_VALID[2]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\OVERFLOW_VALID[1]_i_1_n_0 ),
        .Q(OVERFLOW_VALID__0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \OVERFLOW_VALID_reg[2] 
       (.C(clk_i),
        .CE(\OVERFLOW_VALID[2]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\OVERFLOW_VALID[2]_i_2_n_0 ),
        .Q(OVERFLOW_VALID__0[2]));
  (* srl_bus_name = "\activity_blocks " *) 
  (* srl_name = "\activity_blocks[0].dutH/PAUSEVAL_DEL1_reg_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    PAUSEVAL_DEL1_reg_srl2
       (.A0(1'b1),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b0),
        .CE(1'b1),
        .CLK(clk_i),
        .D(FC_TRANS_PAUSEVAL),
        .Q(PAUSEVAL_DEL1_reg_srl2_n_0));
  FDRE #(
    .INIT(1'b0)) 
    PAUSEVAL_DEL2_reg__0
       (.C(clk_i),
        .CE(1'b1),
        .D(PAUSEVAL_DEL1_reg_srl2_n_0),
        .Q(PAUSEVAL_DEL2),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[0] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[0]),
        .Q(TXC[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[1] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[1]),
        .Q(TXC[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[2] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[2]),
        .Q(TXC[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[3] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[3]),
        .Q(TXC[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[4] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[4]),
        .Q(TXC[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[5] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[5]),
        .Q(TXC[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[6] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[6]),
        .Q(TXC[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXC_reg[7] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_VALID_DEL15[7]),
        .Q(TXC[7]),
        .R(1'b0));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL1_reg[60] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(1'b1),
        .Q(TXD_PAUSE_DEL1));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[0] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[0]),
        .Q(TXD_PAUSE_DEL2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[10] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[10]),
        .Q(TXD_PAUSE_DEL2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[11] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[11]),
        .Q(TXD_PAUSE_DEL2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[12] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[12]),
        .Q(TXD_PAUSE_DEL2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[13] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[13]),
        .Q(TXD_PAUSE_DEL2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[14] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[14]),
        .Q(TXD_PAUSE_DEL2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[15] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[15]),
        .Q(TXD_PAUSE_DEL2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[1] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[1]),
        .Q(TXD_PAUSE_DEL2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[2] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[2]),
        .Q(TXD_PAUSE_DEL2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[3] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[3]),
        .Q(TXD_PAUSE_DEL2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[4] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[4]),
        .Q(TXD_PAUSE_DEL2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[5] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[5]),
        .Q(TXD_PAUSE_DEL2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[6] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[6]),
        .Q(TXD_PAUSE_DEL2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[7] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[7]),
        .Q(TXD_PAUSE_DEL2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[8] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[8]),
        .Q(TXD_PAUSE_DEL2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \TXD_PAUSE_DEL2_reg[9] 
       (.C(clk_i),
        .CE(FC_TRANS_PAUSEVAL),
        .CLR(rst_i),
        .D(FC_TRANS_PAUSEDATA[9]),
        .Q(TXD_PAUSE_DEL2[9]));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[0] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[0]),
        .Q(TXD[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[10] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[10]),
        .Q(TXD[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[11] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[11]),
        .Q(TXD[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[12] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[12]),
        .Q(TXD[12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[13] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[13]),
        .Q(TXD[13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[14] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[14]),
        .Q(TXD[14]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[15] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[15]),
        .Q(TXD[15]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[16] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[16]),
        .Q(TXD[16]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[17] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[17]),
        .Q(TXD[17]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[18] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[18]),
        .Q(TXD[18]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[19] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[19]),
        .Q(TXD[19]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[1] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[1]),
        .Q(TXD[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[20] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[20]),
        .Q(TXD[20]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[21] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[21]),
        .Q(TXD[21]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[22] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[22]),
        .Q(TXD[22]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[23] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[23]),
        .Q(TXD[23]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[24] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[24]),
        .Q(TXD[24]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[25] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[25]),
        .Q(TXD[25]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[26] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[26]),
        .Q(TXD[26]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[27] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[27]),
        .Q(TXD[27]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[28] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[28]),
        .Q(TXD[28]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[29] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[29]),
        .Q(TXD[29]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[2] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[2]),
        .Q(TXD[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[30] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[30]),
        .Q(TXD[30]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[31] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[31]),
        .Q(TXD[31]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[32] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[32]),
        .Q(TXD[32]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[33] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[33]),
        .Q(TXD[33]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[34] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[34]),
        .Q(TXD[34]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[35] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[35]),
        .Q(TXD[35]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[36] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[36]),
        .Q(TXD[36]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[37] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[37]),
        .Q(TXD[37]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[38] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[38]),
        .Q(TXD[38]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[39] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[39]),
        .Q(TXD[39]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[3] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[3]),
        .Q(TXD[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[40] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[40]),
        .Q(TXD[40]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[41] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[41]),
        .Q(TXD[41]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[42] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[42]),
        .Q(TXD[42]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[43] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[43]),
        .Q(TXD[43]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[44] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[44]),
        .Q(TXD[44]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[45] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[45]),
        .Q(TXD[45]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[46] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[46]),
        .Q(TXD[46]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[47] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[47]),
        .Q(TXD[47]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[48] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[48]),
        .Q(TXD[48]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[49] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[49]),
        .Q(TXD[49]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[4] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[4]),
        .Q(TXD[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[50] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[50]),
        .Q(TXD[50]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[51] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[51]),
        .Q(TXD[51]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[52] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[52]),
        .Q(TXD[52]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[53] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[53]),
        .Q(TXD[53]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[54] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[54]),
        .Q(TXD[54]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[55] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[55]),
        .Q(TXD[55]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[56] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[56]),
        .Q(TXD[56]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[57] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[57]),
        .Q(TXD[57]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[58] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[58]),
        .Q(TXD[58]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[59] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[59]),
        .Q(TXD[59]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[5] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[5]),
        .Q(TXD[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[60] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[60]),
        .Q(TXD[60]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[61] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[61]),
        .Q(TXD[61]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[62] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[62]),
        .Q(TXD[62]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[63] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[63]),
        .Q(TXD[63]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[6] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[6]),
        .Q(TXD[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[7] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[7]),
        .Q(TXD[7]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[8] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[8]),
        .Q(TXD[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXD_reg[9] 
       (.C(clk_i),
        .CE(E),
        .D(TX_DATA_DEL15[9]),
        .Q(TXD[9]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(1'b0),
        .Q(TXSTATREGPLUS[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[10] ),
        .Q(TXSTATREGPLUS[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[11] ),
        .Q(TXSTATREGPLUS[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[12] ),
        .Q(TXSTATREGPLUS[12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[13] ),
        .Q(TXSTATREGPLUS[13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[14] ),
        .Q(TXSTATREGPLUS[14]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[15] ),
        .Q(TXSTATREGPLUS[15]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[16] ),
        .Q(TXSTATREGPLUS[16]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[17] ),
        .Q(TXSTATREGPLUS[17]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[18] ),
        .Q(TXSTATREGPLUS[18]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[19] ),
        .Q(TXSTATREGPLUS[19]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[1] ),
        .Q(TXSTATREGPLUS[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(1'b0),
        .Q(TXSTATREGPLUS[20]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(1'b0),
        .Q(TXSTATREGPLUS[21]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(1'b0),
        .Q(TXSTATREGPLUS[22]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(1'b0),
        .Q(TXSTATREGPLUS[23]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[24] ),
        .Q(TXSTATREGPLUS[24]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[2] ),
        .Q(TXSTATREGPLUS[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[3] ),
        .Q(TXSTATREGPLUS[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[4] ),
        .Q(TXSTATREGPLUS[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[5] ),
        .Q(TXSTATREGPLUS[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[6] ),
        .Q(TXSTATREGPLUS[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[7] ),
        .Q(TXSTATREGPLUS[7]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[8] ),
        .Q(TXSTATREGPLUS[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TXSTATREGPLUS_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\txstatplus_int_reg_n_0_[9] ),
        .Q(TXSTATREGPLUS[9]),
        .R(1'b0));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[0]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[0]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[0]),
        .Q(\TX_DATA_DEL11_reg[0]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[10]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[10]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[10]),
        .Q(\TX_DATA_DEL11_reg[10]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[11]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[11]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[11]),
        .Q(\TX_DATA_DEL11_reg[11]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[12]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[12]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[12]),
        .Q(\TX_DATA_DEL11_reg[12]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[13]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[13]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[13]),
        .Q(\TX_DATA_DEL11_reg[13]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[14]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[14]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[14]),
        .Q(\TX_DATA_DEL11_reg[14]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[15]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[15]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[15]),
        .Q(\TX_DATA_DEL11_reg[15]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[16]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[16]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[16]),
        .Q(\TX_DATA_DEL11_reg[16]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[17]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[17]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[17]),
        .Q(\TX_DATA_DEL11_reg[17]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[18]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[18]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[18]),
        .Q(\TX_DATA_DEL11_reg[18]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[19]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[19]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[19]),
        .Q(\TX_DATA_DEL11_reg[19]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[1]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[1]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[1]),
        .Q(\TX_DATA_DEL11_reg[1]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[20]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[20]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[20]),
        .Q(\TX_DATA_DEL11_reg[20]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[21]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[21]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[21]),
        .Q(\TX_DATA_DEL11_reg[21]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[22]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[22]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[22]),
        .Q(\TX_DATA_DEL11_reg[22]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[23]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[23]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[23]),
        .Q(\TX_DATA_DEL11_reg[23]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[24]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[24]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[24]),
        .Q(\TX_DATA_DEL11_reg[24]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[25]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[25]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[25]),
        .Q(\TX_DATA_DEL11_reg[25]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[26]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[26]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[26]),
        .Q(\TX_DATA_DEL11_reg[26]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[27]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[27]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[27]),
        .Q(\TX_DATA_DEL11_reg[27]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[28]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[28]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[28]),
        .Q(\TX_DATA_DEL11_reg[28]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[29]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[29]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[29]),
        .Q(\TX_DATA_DEL11_reg[29]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[2]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[2]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[2]),
        .Q(\TX_DATA_DEL11_reg[2]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[30]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[30]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[30]),
        .Q(\TX_DATA_DEL11_reg[30]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[31]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[31]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[31]),
        .Q(\TX_DATA_DEL11_reg[31]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[32]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[32]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[32]),
        .Q(\TX_DATA_DEL11_reg[32]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[33]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[33]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[33]),
        .Q(\TX_DATA_DEL11_reg[33]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[34]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[34]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[34]),
        .Q(\TX_DATA_DEL11_reg[34]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[35]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[35]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[35]),
        .Q(\TX_DATA_DEL11_reg[35]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[36]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[36]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[36]),
        .Q(\TX_DATA_DEL11_reg[36]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[37]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[37]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[37]),
        .Q(\TX_DATA_DEL11_reg[37]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[38]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[38]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[38]),
        .Q(\TX_DATA_DEL11_reg[38]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[39]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[39]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[39]),
        .Q(\TX_DATA_DEL11_reg[39]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[3]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[3]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[3]),
        .Q(\TX_DATA_DEL11_reg[3]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[40]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[40]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[40]),
        .Q(\TX_DATA_DEL11_reg[40]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[41]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[41]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[41]),
        .Q(\TX_DATA_DEL11_reg[41]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[42]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[42]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[42]),
        .Q(\TX_DATA_DEL11_reg[42]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[43]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[43]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[43]),
        .Q(\TX_DATA_DEL11_reg[43]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[44]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[44]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[44]),
        .Q(\TX_DATA_DEL11_reg[44]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[45]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[45]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[45]),
        .Q(\TX_DATA_DEL11_reg[45]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[46]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[46]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[46]),
        .Q(\TX_DATA_DEL11_reg[46]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[47]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[47]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[47]),
        .Q(\TX_DATA_DEL11_reg[47]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[48]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[48]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[48]),
        .Q(\TX_DATA_DEL11_reg[48]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[49]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[49]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[49]),
        .Q(\TX_DATA_DEL11_reg[49]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[4]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[4]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[4]),
        .Q(\TX_DATA_DEL11_reg[4]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[50]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[50]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[50]),
        .Q(\TX_DATA_DEL11_reg[50]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[51]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[51]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[51]),
        .Q(\TX_DATA_DEL11_reg[51]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[52]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[52]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[52]),
        .Q(\TX_DATA_DEL11_reg[52]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[53]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[53]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[53]),
        .Q(\TX_DATA_DEL11_reg[53]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[54]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[54]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[54]),
        .Q(\TX_DATA_DEL11_reg[54]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[55]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[55]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[55]),
        .Q(\TX_DATA_DEL11_reg[55]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[56]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[56]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[56]),
        .Q(\TX_DATA_DEL11_reg[56]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[57]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[57]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[57]),
        .Q(\TX_DATA_DEL11_reg[57]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[58]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[58]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[58]),
        .Q(\TX_DATA_DEL11_reg[58]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[59]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[59]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[59]),
        .Q(\TX_DATA_DEL11_reg[59]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[5]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[5]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[5]),
        .Q(\TX_DATA_DEL11_reg[5]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[60]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[60]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[60]),
        .Q(\TX_DATA_DEL11_reg[60]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[61]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[61]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[61]),
        .Q(\TX_DATA_DEL11_reg[61]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[62]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[62]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[62]),
        .Q(\TX_DATA_DEL11_reg[62]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[63]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[63]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[63]),
        .Q(\TX_DATA_DEL11_reg[63]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[6]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[6]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[6]),
        .Q(\TX_DATA_DEL11_reg[6]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[7]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[7]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[7]),
        .Q(\TX_DATA_DEL11_reg[7]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[8]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[8]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[8]),
        .Q(\TX_DATA_DEL11_reg[8]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_DEL11_reg[9]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_DEL11_reg[9]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_DEL2[9]),
        .Q(\TX_DATA_DEL11_reg[9]_srl9_activity_blocks_c_7_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[0]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[0]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[0]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[10]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[10]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[10]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[11]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[11]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[11]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[12]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[12]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[12]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[13]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[13]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[13]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[14]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[14]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[14]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[15]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[15]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[15]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[16]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[16]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[16]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[17]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[17]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[17]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[18]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[18]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[18]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[19]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[19]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[19]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[1]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[1]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[1]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[20]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[20]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[20]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[21]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[21]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[21]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[22]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[22]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[22]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[23]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[23]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[23]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[24]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[24]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[24]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[25]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[25]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[25]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[26]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[26]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[26]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[27]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[27]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[27]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[28]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[28]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[28]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[29]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[29]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[29]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[2]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[2]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[2]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[30]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[30]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[30]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[31]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[31]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[31]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[32]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[32]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[32]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[33]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[33]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[33]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[34]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[34]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[34]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[35]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[35]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[35]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[36]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[36]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[36]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[37]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[37]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[37]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[38]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[38]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[38]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[39]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[39]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[39]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[3]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[3]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[3]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[40]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[40]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[40]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[41]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[41]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[41]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[42]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[42]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[42]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[43]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[43]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[43]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[44]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[44]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[44]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[45]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[45]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[45]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[46]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[46]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[46]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[47]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[47]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[47]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[48]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[48]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[48]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[49]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[49]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[49]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[4]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[4]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[4]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[50]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[50]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[50]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[51]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[51]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[51]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[52]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[52]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[52]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[53]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[53]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[53]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[54]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[54]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[54]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[55]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[55]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[55]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[56]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[56]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[56]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[57]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[57]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[57]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[58]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[58]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[58]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[59]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[59]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[59]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[5]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[5]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[5]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[60]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[60]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[60]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[61]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[61]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[61]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[62]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[62]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[62]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[63]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[63]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[63]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[6]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[6]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[6]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[7]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[7]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[7]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[8]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[8]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[8]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL12_reg[9]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_DEL11_reg[9]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_DEL12_reg[9]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__71_n_0),
        .Q(TX_DATA_DEL13[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__61_n_0),
        .Q(TX_DATA_DEL13[10]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__60_n_0),
        .Q(TX_DATA_DEL13[11]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__59_n_0),
        .Q(TX_DATA_DEL13[12]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__58_n_0),
        .Q(TX_DATA_DEL13[13]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__57_n_0),
        .Q(TX_DATA_DEL13[14]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__56_n_0),
        .Q(TX_DATA_DEL13[15]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__55_n_0),
        .Q(TX_DATA_DEL13[16]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__54_n_0),
        .Q(TX_DATA_DEL13[17]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__53_n_0),
        .Q(TX_DATA_DEL13[18]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__52_n_0),
        .Q(TX_DATA_DEL13[19]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__70_n_0),
        .Q(TX_DATA_DEL13[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__51_n_0),
        .Q(TX_DATA_DEL13[20]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__50_n_0),
        .Q(TX_DATA_DEL13[21]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__49_n_0),
        .Q(TX_DATA_DEL13[22]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__48_n_0),
        .Q(TX_DATA_DEL13[23]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__47_n_0),
        .Q(TX_DATA_DEL13[24]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__46_n_0),
        .Q(TX_DATA_DEL13[25]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__45_n_0),
        .Q(TX_DATA_DEL13[26]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__44_n_0),
        .Q(TX_DATA_DEL13[27]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__43_n_0),
        .Q(TX_DATA_DEL13[28]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__42_n_0),
        .Q(TX_DATA_DEL13[29]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__69_n_0),
        .Q(TX_DATA_DEL13[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__41_n_0),
        .Q(TX_DATA_DEL13[30]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__40_n_0),
        .Q(TX_DATA_DEL13[31]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__39_n_0),
        .Q(TX_DATA_DEL13[32]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__38_n_0),
        .Q(TX_DATA_DEL13[33]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__37_n_0),
        .Q(TX_DATA_DEL13[34]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__36_n_0),
        .Q(TX_DATA_DEL13[35]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__35_n_0),
        .Q(TX_DATA_DEL13[36]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__34_n_0),
        .Q(TX_DATA_DEL13[37]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__33_n_0),
        .Q(TX_DATA_DEL13[38]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__32_n_0),
        .Q(TX_DATA_DEL13[39]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__68_n_0),
        .Q(TX_DATA_DEL13[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__31_n_0),
        .Q(TX_DATA_DEL13[40]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__30_n_0),
        .Q(TX_DATA_DEL13[41]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__29_n_0),
        .Q(TX_DATA_DEL13[42]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__28_n_0),
        .Q(TX_DATA_DEL13[43]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__27_n_0),
        .Q(TX_DATA_DEL13[44]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__26_n_0),
        .Q(TX_DATA_DEL13[45]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__25_n_0),
        .Q(TX_DATA_DEL13[46]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__24_n_0),
        .Q(TX_DATA_DEL13[47]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__23_n_0),
        .Q(TX_DATA_DEL13[48]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__22_n_0),
        .Q(TX_DATA_DEL13[49]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__67_n_0),
        .Q(TX_DATA_DEL13[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__21_n_0),
        .Q(TX_DATA_DEL13[50]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__20_n_0),
        .Q(TX_DATA_DEL13[51]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__19_n_0),
        .Q(TX_DATA_DEL13[52]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__18_n_0),
        .Q(TX_DATA_DEL13[53]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__17_n_0),
        .Q(TX_DATA_DEL13[54]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__16_n_0),
        .Q(TX_DATA_DEL13[55]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__15_n_0),
        .Q(TX_DATA_DEL13[56]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__14_n_0),
        .Q(TX_DATA_DEL13[57]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__13_n_0),
        .Q(TX_DATA_DEL13[58]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__12_n_0),
        .Q(TX_DATA_DEL13[59]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__66_n_0),
        .Q(TX_DATA_DEL13[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__11_n_0),
        .Q(TX_DATA_DEL13[60]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__10_n_0),
        .Q(TX_DATA_DEL13[61]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__9_n_0),
        .Q(TX_DATA_DEL13[62]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__8_n_0),
        .Q(TX_DATA_DEL13[63]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__65_n_0),
        .Q(TX_DATA_DEL13[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__64_n_0),
        .Q(TX_DATA_DEL13[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__63_n_0),
        .Q(TX_DATA_DEL13[8]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL13_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__62_n_0),
        .Q(TX_DATA_DEL13[9]));
  (* SOFT_HLUTNM = "soft_lutpair442" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    \TX_DATA_DEL14[15]_i_2 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[58]_i_3_n_0 ),
        .I2(\TX_DATA_DEL14[50]_i_3_n_0 ),
        .I3(\TX_DATA_DEL14[63]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[18]_i_4 
       (.I0(\OVERFLOW_DATA_reg_n_0_[18] ),
        .I1(append_end_frame),
        .I2(TX_DATA_DEL13[18]),
        .O(\TX_DATA_DEL14[18]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair442" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \TX_DATA_DEL14[23]_i_2 
       (.I0(\TX_DATA_DEL14[50]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[58]_i_3_n_0 ),
        .I2(TX_DATA_VALID_DEL13),
        .O(\TX_DATA_DEL14[23]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair487" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[25]_i_4 
       (.I0(\OVERFLOW_DATA_reg_n_0_[25] ),
        .I1(append_end_frame),
        .I2(TX_DATA_DEL13[25]),
        .O(\TX_DATA_DEL14[25]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair488" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \TX_DATA_DEL14[33]_i_4 
       (.I0(\OVERFLOW_DATA_reg_n_0_[33] ),
        .I1(append_end_frame),
        .I2(TX_DATA_DEL13[33]),
        .O(\TX_DATA_DEL14[33]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair447" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[33]_i_6 
       (.I0(fcs_enabled_int),
        .I1(txstatplus_int),
        .O(\TX_DATA_DEL14[33]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair488" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \TX_DATA_DEL14[39]_i_3 
       (.I0(txstatplus_int0_out[1]),
        .I1(\OVERFLOW_DATA_reg_n_0_[39] ),
        .I2(append_end_frame),
        .O(\TX_DATA_DEL14[39]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5555555544545555)) 
    \TX_DATA_DEL14[39]_i_5 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(\TX_DATA_DEL14[63]_i_8_n_0 ),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[2]),
        .I5(TX_DATA_VALID_DEL13__0[6]),
        .O(\TX_DATA_DEL14[39]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h4100FFFF)) 
    \TX_DATA_DEL14[41]_i_5 
       (.I0(TX_DATA_VALID_DEL13__0[6]),
        .I1(TX_DATA_VALID_DEL13__0[5]),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .I3(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .I4(TX_DATA_DEL13[41]),
        .O(\TX_DATA_DEL14[41]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \TX_DATA_DEL14[47]_i_3 
       (.I0(\TX_DATA_DEL14[58]_i_3_n_0 ),
        .I1(\TX_DATA_DEL14[50]_i_3_n_0 ),
        .I2(TX_DATA_DEL13[47]),
        .O(\TX_DATA_DEL14[47]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair419" *) 
  LUT5 #(
    .INIT(32'hBAABAAAA)) 
    \TX_DATA_DEL14[48]_i_5 
       (.I0(TX_DATA_DEL13[48]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[48]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FF700004004)) 
    \TX_DATA_DEL14[48]_i_6 
       (.I0(\OVERFLOW_DATA[8]_i_2_n_0 ),
        .I1(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .I3(TX_DATA_VALID_DEL13__0[5]),
        .I4(TX_DATA_VALID_DEL13__0[6]),
        .I5(TX_DATA_DEL13[48]),
        .O(\TX_DATA_DEL14[48]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBAABAAAA)) 
    \TX_DATA_DEL14[49]_i_5 
       (.I0(TX_DATA_DEL13[49]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[49]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2AA2AAAAEAAE)) 
    \TX_DATA_DEL14[49]_i_6 
       (.I0(TX_DATA_DEL13[49]),
        .I1(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .I3(TX_DATA_VALID_DEL13__0[5]),
        .I4(TX_DATA_VALID_DEL13__0[6]),
        .I5(\TX_DATA_DEL14[33]_i_6_n_0 ),
        .O(\TX_DATA_DEL14[49]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair419" *) 
  LUT4 #(
    .INIT(16'h0082)) 
    \TX_DATA_DEL14[50]_i_3 
       (.I0(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[4]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .O(\TX_DATA_DEL14[50]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair427" *) 
  LUT5 #(
    .INIT(32'h80800009)) 
    \TX_DATA_DEL14[50]_i_5 
       (.I0(TX_DATA_VALID_DEL13__0[0]),
        .I1(TX_DATA_VALID_DEL13__0[1]),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[2]),
        .O(\TX_DATA_DEL14[50]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h8AA8AAAA)) 
    \TX_DATA_DEL14[51]_i_5 
       (.I0(TX_DATA_DEL13[51]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[51]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair443" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \TX_DATA_DEL14[52]_i_3 
       (.I0(fcs_enabled_int),
        .I1(\TX_DATA_DEL14[63]_i_5_n_0 ),
        .I2(\TX_DATA_DEL14[50]_i_3_n_0 ),
        .I3(TX_DATA_DEL13[52]),
        .O(\TX_DATA_DEL14[52]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair444" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \TX_DATA_DEL14[53]_i_3 
       (.I0(fcs_enabled_int),
        .I1(\TX_DATA_DEL14[63]_i_5_n_0 ),
        .I2(\TX_DATA_DEL14[50]_i_3_n_0 ),
        .I3(TX_DATA_DEL13[53]),
        .O(\TX_DATA_DEL14[53]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair423" *) 
  LUT5 #(
    .INIT(32'hDFFDFFFF)) 
    \TX_DATA_DEL14[54]_i_5 
       (.I0(fcs_enabled_int),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[54]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h8AA8AAAA)) 
    \TX_DATA_DEL14[54]_i_6 
       (.I0(TX_DATA_DEL13[54]),
        .I1(TX_DATA_VALID_DEL13__0[6]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[54]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair443" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \TX_DATA_DEL14[55]_i_3 
       (.I0(fcs_enabled_int),
        .I1(\TX_DATA_DEL14[63]_i_5_n_0 ),
        .I2(\TX_DATA_DEL14[50]_i_3_n_0 ),
        .I3(TX_DATA_DEL13[55]),
        .O(\TX_DATA_DEL14[55]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000A800FCFCA8FC)) 
    \TX_DATA_DEL14[57]_i_6 
       (.I0(\OVERFLOW_DATA[8]_i_2_n_0 ),
        .I1(\TX_DATA_VALID_DEL14[6]_i_3_n_0 ),
        .I2(\TX_DATA_DEL14[57]_i_8_n_0 ),
        .I3(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .I4(\TX_DATA_DEL14[57]_i_7_n_0 ),
        .I5(TX_DATA_DEL13[57]),
        .O(\TX_DATA_DEL14[57]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair420" *) 
  LUT3 #(
    .INIT(8'hBE)) 
    \TX_DATA_DEL14[57]_i_7 
       (.I0(TX_DATA_VALID_DEL13__0[6]),
        .I1(TX_DATA_VALID_DEL13__0[5]),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .O(\TX_DATA_DEL14[57]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair422" *) 
  LUT5 #(
    .INIT(32'h7FFFFFF2)) 
    \TX_DATA_DEL14[57]_i_8 
       (.I0(TX_DATA_VALID_DEL13__0[3]),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(TX_DATA_VALID_DEL13__0[6]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[5]),
        .O(\TX_DATA_DEL14[57]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4400040400000000)) 
    \TX_DATA_DEL14[58]_i_3 
       (.I0(TX_DATA_VALID_DEL13__0[6]),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .I5(\TX_DATA_DEL14[58]_i_7_n_0 ),
        .O(\TX_DATA_DEL14[58]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair425" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[58]_i_5 
       (.I0(txstatplus_int0_out[1]),
        .I1(TX_DATA_VALID_DEL13),
        .O(\TX_DATA_DEL14[58]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair430" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \TX_DATA_DEL14[58]_i_6 
       (.I0(append_end_frame),
        .I1(txstatplus_int0_out[1]),
        .O(\TX_DATA_DEL14[58]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_DEL14[58]_i_7 
       (.I0(TX_DATA_VALID_DEL13__0[1]),
        .I1(TX_DATA_VALID_DEL13__0[0]),
        .O(\TX_DATA_DEL14[58]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000510000000000)) 
    \TX_DATA_DEL14[63]_i_4 
       (.I0(\TX_DATA_DEL14[63]_i_8_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[5]),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(TX_DATA_VALID_DEL13__0[6]),
        .I5(\TX_DATA_DEL14[58]_i_5_n_0 ),
        .O(\TX_DATA_DEL14[63]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4001000000010001)) 
    \TX_DATA_DEL14[63]_i_5 
       (.I0(\TX_DATA_VALID_DEL14[6]_i_3_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[5]),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .I4(TX_DATA_VALID_DEL13__0[2]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(\TX_DATA_DEL14[63]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88A8AAAA)) 
    \TX_DATA_DEL14[63]_i_7 
       (.I0(\TX_DATA_DEL14[58]_i_5_n_0 ),
        .I1(\TX_DATA_DEL14[63]_i_8_n_0 ),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(TX_DATA_VALID_DEL13__0[2]),
        .I5(TX_DATA_VALID_DEL13__0[6]),
        .O(\TX_DATA_DEL14[63]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair427" *) 
  LUT4 #(
    .INIT(16'h77F7)) 
    \TX_DATA_DEL14[63]_i_8 
       (.I0(TX_DATA_VALID_DEL13__0[0]),
        .I1(TX_DATA_VALID_DEL13__0[1]),
        .I2(TX_DATA_VALID_DEL13__0[4]),
        .I3(TX_DATA_VALID_DEL13__0[3]),
        .O(\TX_DATA_DEL14[63]_i_8_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_88),
        .Q(\TX_DATA_DEL14_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_78),
        .Q(\TX_DATA_DEL14_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_77),
        .Q(\TX_DATA_DEL14_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_76),
        .Q(\TX_DATA_DEL14_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_75),
        .Q(\TX_DATA_DEL14_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_74),
        .Q(\TX_DATA_DEL14_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_73),
        .Q(\TX_DATA_DEL14_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_72),
        .Q(\TX_DATA_DEL14_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_71),
        .Q(\TX_DATA_DEL14_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_70),
        .Q(\TX_DATA_DEL14_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_69),
        .Q(\TX_DATA_DEL14_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_87),
        .Q(\TX_DATA_DEL14_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_68),
        .Q(\TX_DATA_DEL14_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_67),
        .Q(\TX_DATA_DEL14_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_66),
        .Q(\TX_DATA_DEL14_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_65),
        .Q(\TX_DATA_DEL14_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_64),
        .Q(\TX_DATA_DEL14_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_63),
        .Q(\TX_DATA_DEL14_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_62),
        .Q(\TX_DATA_DEL14_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_61),
        .Q(\TX_DATA_DEL14_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_60),
        .Q(\TX_DATA_DEL14_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_59),
        .Q(\TX_DATA_DEL14_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_86),
        .Q(\TX_DATA_DEL14_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_58),
        .Q(\TX_DATA_DEL14_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_57),
        .Q(\TX_DATA_DEL14_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_56),
        .Q(\TX_DATA_DEL14_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_55),
        .Q(\TX_DATA_DEL14_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_54),
        .Q(\TX_DATA_DEL14_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_53),
        .Q(\TX_DATA_DEL14_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_52),
        .Q(\TX_DATA_DEL14_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_51),
        .Q(\TX_DATA_DEL14_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_50),
        .Q(\TX_DATA_DEL14_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_49),
        .Q(\TX_DATA_DEL14_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_85),
        .Q(\TX_DATA_DEL14_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_48),
        .Q(\TX_DATA_DEL14_reg_n_0_[40] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_47),
        .Q(\TX_DATA_DEL14_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_46),
        .Q(\TX_DATA_DEL14_reg_n_0_[42] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_45),
        .Q(\TX_DATA_DEL14_reg_n_0_[43] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_44),
        .Q(\TX_DATA_DEL14_reg_n_0_[44] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_43),
        .Q(\TX_DATA_DEL14_reg_n_0_[45] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_42),
        .Q(\TX_DATA_DEL14_reg_n_0_[46] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_41),
        .Q(\TX_DATA_DEL14_reg_n_0_[47] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_40),
        .Q(\TX_DATA_DEL14_reg_n_0_[48] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_39),
        .Q(\TX_DATA_DEL14_reg_n_0_[49] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_84),
        .Q(\TX_DATA_DEL14_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_38),
        .Q(\TX_DATA_DEL14_reg_n_0_[50] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_37),
        .Q(\TX_DATA_DEL14_reg_n_0_[51] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_36),
        .Q(\TX_DATA_DEL14_reg_n_0_[52] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_35),
        .Q(\TX_DATA_DEL14_reg_n_0_[53] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_34),
        .Q(\TX_DATA_DEL14_reg_n_0_[54] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_33),
        .Q(\TX_DATA_DEL14_reg_n_0_[55] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_32),
        .Q(\TX_DATA_DEL14_reg_n_0_[56] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_31),
        .Q(\TX_DATA_DEL14_reg_n_0_[57] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_30),
        .Q(\TX_DATA_DEL14_reg_n_0_[58] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_29),
        .Q(\TX_DATA_DEL14_reg_n_0_[59] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_83),
        .Q(\TX_DATA_DEL14_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_28),
        .Q(\TX_DATA_DEL14_reg_n_0_[60] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_27),
        .Q(\TX_DATA_DEL14_reg_n_0_[61] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_26),
        .Q(\TX_DATA_DEL14_reg_n_0_[62] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_25),
        .Q(\TX_DATA_DEL14_reg_n_0_[63] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_82),
        .Q(\TX_DATA_DEL14_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_81),
        .Q(\TX_DATA_DEL14_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_80),
        .Q(\TX_DATA_DEL14_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL14_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_CRC8_n_79),
        .Q(\TX_DATA_DEL14_reg_n_0_[9] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[0] ),
        .Q(TX_DATA_DEL15[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[10] ),
        .Q(TX_DATA_DEL15[10]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[11] ),
        .Q(TX_DATA_DEL15[11]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[12] ),
        .Q(TX_DATA_DEL15[12]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[13] ),
        .Q(TX_DATA_DEL15[13]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[14] ),
        .Q(TX_DATA_DEL15[14]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[15] ),
        .Q(TX_DATA_DEL15[15]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[16] ),
        .Q(TX_DATA_DEL15[16]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[17] ),
        .Q(TX_DATA_DEL15[17]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[18] ),
        .Q(TX_DATA_DEL15[18]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[19] ),
        .Q(TX_DATA_DEL15[19]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[1] ),
        .Q(TX_DATA_DEL15[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[20] ),
        .Q(TX_DATA_DEL15[20]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[21] ),
        .Q(TX_DATA_DEL15[21]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[22] ),
        .Q(TX_DATA_DEL15[22]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[23] ),
        .Q(TX_DATA_DEL15[23]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[24] ),
        .Q(TX_DATA_DEL15[24]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[25] ),
        .Q(TX_DATA_DEL15[25]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[26] ),
        .Q(TX_DATA_DEL15[26]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[27] ),
        .Q(TX_DATA_DEL15[27]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[28] ),
        .Q(TX_DATA_DEL15[28]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[29] ),
        .Q(TX_DATA_DEL15[29]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[2] ),
        .Q(TX_DATA_DEL15[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[30] ),
        .Q(TX_DATA_DEL15[30]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[31] ),
        .Q(TX_DATA_DEL15[31]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[32] ),
        .Q(TX_DATA_DEL15[32]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[33] ),
        .Q(TX_DATA_DEL15[33]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[34] ),
        .Q(TX_DATA_DEL15[34]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[35] ),
        .Q(TX_DATA_DEL15[35]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[36] ),
        .Q(TX_DATA_DEL15[36]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[37] ),
        .Q(TX_DATA_DEL15[37]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[38] ),
        .Q(TX_DATA_DEL15[38]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[39] ),
        .Q(TX_DATA_DEL15[39]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[3] ),
        .Q(TX_DATA_DEL15[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[40] ),
        .Q(TX_DATA_DEL15[40]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[41] ),
        .Q(TX_DATA_DEL15[41]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[42] ),
        .Q(TX_DATA_DEL15[42]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[43] ),
        .Q(TX_DATA_DEL15[43]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[44] ),
        .Q(TX_DATA_DEL15[44]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[45] ),
        .Q(TX_DATA_DEL15[45]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[46] ),
        .Q(TX_DATA_DEL15[46]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[47] ),
        .Q(TX_DATA_DEL15[47]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[48] ),
        .Q(TX_DATA_DEL15[48]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[49] ),
        .Q(TX_DATA_DEL15[49]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[4] ),
        .Q(TX_DATA_DEL15[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[50] ),
        .Q(TX_DATA_DEL15[50]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[51] ),
        .Q(TX_DATA_DEL15[51]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[52] ),
        .Q(TX_DATA_DEL15[52]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[53] ),
        .Q(TX_DATA_DEL15[53]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[54] ),
        .Q(TX_DATA_DEL15[54]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[55] ),
        .Q(TX_DATA_DEL15[55]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[56] ),
        .Q(TX_DATA_DEL15[56]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[57] ),
        .Q(TX_DATA_DEL15[57]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[58] ),
        .Q(TX_DATA_DEL15[58]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[59] ),
        .Q(TX_DATA_DEL15[59]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[5] ),
        .Q(TX_DATA_DEL15[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[60] ),
        .Q(TX_DATA_DEL15[60]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[61] ),
        .Q(TX_DATA_DEL15[61]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[62] ),
        .Q(TX_DATA_DEL15[62]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[63] ),
        .Q(TX_DATA_DEL15[63]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[6] ),
        .Q(TX_DATA_DEL15[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[7] ),
        .Q(TX_DATA_DEL15[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[8] ),
        .Q(TX_DATA_DEL15[8]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL15_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_DEL14_reg_n_0_[9] ),
        .Q(TX_DATA_DEL15[9]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[0] ),
        .Q(TX_DATA_DEL1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[10] ),
        .Q(TX_DATA_DEL1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[11] ),
        .Q(TX_DATA_DEL1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[12] ),
        .Q(TX_DATA_DEL1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[13] ),
        .Q(TX_DATA_DEL1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[14] ),
        .Q(TX_DATA_DEL1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[15] ),
        .Q(TX_DATA_DEL1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[16] ),
        .Q(TX_DATA_DEL1[16]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[17] ),
        .Q(TX_DATA_DEL1[17]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[18] ),
        .Q(TX_DATA_DEL1[18]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[19] ),
        .Q(TX_DATA_DEL1[19]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[1] ),
        .Q(TX_DATA_DEL1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[20] ),
        .Q(TX_DATA_DEL1[20]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[21] ),
        .Q(TX_DATA_DEL1[21]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[22] ),
        .Q(TX_DATA_DEL1[22]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[23] ),
        .Q(TX_DATA_DEL1[23]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[24] ),
        .Q(TX_DATA_DEL1[24]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[25] ),
        .Q(TX_DATA_DEL1[25]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[26] ),
        .Q(TX_DATA_DEL1[26]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[27] ),
        .Q(TX_DATA_DEL1[27]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[28] ),
        .Q(TX_DATA_DEL1[28]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[29] ),
        .Q(TX_DATA_DEL1[29]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[2] ),
        .Q(TX_DATA_DEL1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[30] ),
        .Q(TX_DATA_DEL1[30]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[31] ),
        .Q(TX_DATA_DEL1[31]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[32] ),
        .Q(TX_DATA_DEL1[32]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[33] ),
        .Q(TX_DATA_DEL1[33]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[34] ),
        .Q(TX_DATA_DEL1[34]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[35] ),
        .Q(TX_DATA_DEL1[35]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[36] ),
        .Q(TX_DATA_DEL1[36]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[37] ),
        .Q(TX_DATA_DEL1[37]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[38] ),
        .Q(TX_DATA_DEL1[38]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[39] ),
        .Q(TX_DATA_DEL1[39]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[3] ),
        .Q(TX_DATA_DEL1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[40] ),
        .Q(TX_DATA_DEL1[40]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[41] ),
        .Q(TX_DATA_DEL1[41]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[42] ),
        .Q(TX_DATA_DEL1[42]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[43] ),
        .Q(TX_DATA_DEL1[43]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[44] ),
        .Q(TX_DATA_DEL1[44]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[45] ),
        .Q(TX_DATA_DEL1[45]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[46] ),
        .Q(TX_DATA_DEL1[46]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[47] ),
        .Q(TX_DATA_DEL1[47]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[48] ),
        .Q(TX_DATA_DEL1[48]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[49] ),
        .Q(TX_DATA_DEL1[49]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[4] ),
        .Q(TX_DATA_DEL1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[50] ),
        .Q(TX_DATA_DEL1[50]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[51] ),
        .Q(TX_DATA_DEL1[51]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[52] ),
        .Q(TX_DATA_DEL1[52]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[53] ),
        .Q(TX_DATA_DEL1[53]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[54] ),
        .Q(TX_DATA_DEL1[54]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[55] ),
        .Q(TX_DATA_DEL1[55]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[56] ),
        .Q(TX_DATA_DEL1[56]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[57] ),
        .Q(TX_DATA_DEL1[57]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[58] ),
        .Q(TX_DATA_DEL1[58]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[59] ),
        .Q(TX_DATA_DEL1[59]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[5] ),
        .Q(TX_DATA_DEL1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[60] ),
        .Q(TX_DATA_DEL1[60]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[61] ),
        .Q(TX_DATA_DEL1[61]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[62] ),
        .Q(TX_DATA_DEL1[62]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[63] ),
        .Q(TX_DATA_DEL1[63]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[6] ),
        .Q(TX_DATA_DEL1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[7] ),
        .Q(TX_DATA_DEL1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[8] ),
        .Q(TX_DATA_DEL1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_REG_reg_n_0_[9] ),
        .Q(TX_DATA_DEL1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[0]),
        .Q(TX_DATA_DEL2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[10]),
        .Q(TX_DATA_DEL2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[11]),
        .Q(TX_DATA_DEL2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[12]),
        .Q(TX_DATA_DEL2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[13]),
        .Q(TX_DATA_DEL2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[14]),
        .Q(TX_DATA_DEL2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[15]),
        .Q(TX_DATA_DEL2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[16]),
        .Q(TX_DATA_DEL2[16]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[17]),
        .Q(TX_DATA_DEL2[17]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[18]),
        .Q(TX_DATA_DEL2[18]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[19]),
        .Q(TX_DATA_DEL2[19]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[1]),
        .Q(TX_DATA_DEL2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[20]),
        .Q(TX_DATA_DEL2[20]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[21]),
        .Q(TX_DATA_DEL2[21]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[22]),
        .Q(TX_DATA_DEL2[22]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[23]),
        .Q(TX_DATA_DEL2[23]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[24]),
        .Q(TX_DATA_DEL2[24]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[25]),
        .Q(TX_DATA_DEL2[25]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[26]),
        .Q(TX_DATA_DEL2[26]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[27]),
        .Q(TX_DATA_DEL2[27]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[28]),
        .Q(TX_DATA_DEL2[28]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[29]),
        .Q(TX_DATA_DEL2[29]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[2]),
        .Q(TX_DATA_DEL2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[30]),
        .Q(TX_DATA_DEL2[30]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[31]),
        .Q(TX_DATA_DEL2[31]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[32]),
        .Q(TX_DATA_DEL2[32]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[33]),
        .Q(TX_DATA_DEL2[33]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[34]),
        .Q(TX_DATA_DEL2[34]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[35]),
        .Q(TX_DATA_DEL2[35]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[36]),
        .Q(TX_DATA_DEL2[36]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[37]),
        .Q(TX_DATA_DEL2[37]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[38]),
        .Q(TX_DATA_DEL2[38]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[39]),
        .Q(TX_DATA_DEL2[39]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[3]),
        .Q(TX_DATA_DEL2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[40]),
        .Q(TX_DATA_DEL2[40]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[41]),
        .Q(TX_DATA_DEL2[41]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[42]),
        .Q(TX_DATA_DEL2[42]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[43]),
        .Q(TX_DATA_DEL2[43]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[44]),
        .Q(TX_DATA_DEL2[44]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[45]),
        .Q(TX_DATA_DEL2[45]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[46]),
        .Q(TX_DATA_DEL2[46]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[47]),
        .Q(TX_DATA_DEL2[47]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[48]),
        .Q(TX_DATA_DEL2[48]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[49]),
        .Q(TX_DATA_DEL2[49]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[4]),
        .Q(TX_DATA_DEL2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[50]),
        .Q(TX_DATA_DEL2[50]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[51]),
        .Q(TX_DATA_DEL2[51]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[52]),
        .Q(TX_DATA_DEL2[52]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[53]),
        .Q(TX_DATA_DEL2[53]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[54]),
        .Q(TX_DATA_DEL2[54]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[55]),
        .Q(TX_DATA_DEL2[55]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[56]),
        .Q(TX_DATA_DEL2[56]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[57]),
        .Q(TX_DATA_DEL2[57]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[58]),
        .Q(TX_DATA_DEL2[58]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[59]),
        .Q(TX_DATA_DEL2[59]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[5]),
        .Q(TX_DATA_DEL2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[60]),
        .Q(TX_DATA_DEL2[60]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[61]),
        .Q(TX_DATA_DEL2[61]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[62]),
        .Q(TX_DATA_DEL2[62]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[63]),
        .Q(TX_DATA_DEL2[63]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[6]),
        .Q(TX_DATA_DEL2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[7]),
        .Q(TX_DATA_DEL2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[8]),
        .Q(TX_DATA_DEL2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_DEL2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_DEL1[9]),
        .Q(TX_DATA_DEL2[9]));
  (* SOFT_HLUTNM = "soft_lutpair431" *) 
  LUT4 #(
    .INIT(16'hB8BB)) 
    \TX_DATA_REG[0]_i_1 
       (.I0(TX_DATA_VALID_DELAY[0]),
        .I1(FRAME_START),
        .I2(shift_pause_data[0]),
        .I3(transmit_pause_frame_valid),
        .O(\TX_DATA_REG[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair432" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \TX_DATA_REG[12]_i_2 
       (.I0(shift_pause_data[12]),
        .I1(transmit_pause_frame_valid),
        .I2(FRAME_START),
        .O(\TX_DATA_REG[12]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair469" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \TX_DATA_REG[14]_i_2 
       (.I0(shift_pause_data[14]),
        .I1(transmit_pause_frame_valid),
        .I2(FRAME_START),
        .O(\TX_DATA_REG[14]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair432" *) 
  LUT4 #(
    .INIT(16'hB8BB)) 
    \TX_DATA_REG[1]_i_1 
       (.I0(TX_DATA_VALID_DELAY[1]),
        .I1(FRAME_START),
        .I2(shift_pause_data[1]),
        .I3(transmit_pause_frame_valid),
        .O(\TX_DATA_REG[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair489" *) 
  LUT3 #(
    .INIT(8'h0D)) 
    \TX_DATA_REG[56]_i_2 
       (.I0(transmit_pause_frame_valid),
        .I1(shift_pause_data[56]),
        .I2(FRAME_START),
        .O(\TX_DATA_REG[56]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair489" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \TX_DATA_REG[60]_i_2 
       (.I0(shift_pause_data[60]),
        .I1(transmit_pause_frame_valid),
        .I2(FRAME_START),
        .O(\TX_DATA_REG[60]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h50110001FFFFFFFF)) 
    \TX_DATA_REG[63]_i_4 
       (.I0(\TX_DATA_REG[63]_i_6_n_0 ),
        .I1(\TX_DATA_VALID_REG_reg_n_0_[7] ),
        .I2(\TX_DATA_VALID_REG_reg_n_0_[5] ),
        .I3(\TX_DATA_VALID_REG_reg_n_0_[6] ),
        .I4(\TX_DATA_VALID_REG_reg_n_0_[4] ),
        .I5(FRAME_START),
        .O(\TX_DATA_REG[63]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair429" *) 
  LUT5 #(
    .INIT(32'h7F77FFF2)) 
    \TX_DATA_REG[63]_i_6 
       (.I0(\TX_DATA_VALID_REG_reg_n_0_[1] ),
        .I1(\TX_DATA_VALID_REG_reg_n_0_[0] ),
        .I2(\TX_DATA_VALID_REG_reg_n_0_[3] ),
        .I3(\TX_DATA_VALID_REG_reg_n_0_[4] ),
        .I4(\TX_DATA_VALID_REG_reg_n_0_[2] ),
        .O(\TX_DATA_REG[63]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair431" *) 
  LUT3 #(
    .INIT(8'h45)) 
    \TX_DATA_REG[9]_i_2 
       (.I0(FRAME_START),
        .I1(shift_pause_data[9]),
        .I2(transmit_pause_frame_valid),
        .O(\TX_DATA_REG[9]_i_2_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[0] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(\TX_DATA_REG[0]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[0] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[10] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_102),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[11] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_101),
        .Q(\TX_DATA_REG_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[12] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_100),
        .Q(\TX_DATA_REG_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[13] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_99),
        .Q(\TX_DATA_REG_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[14] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_98),
        .Q(\TX_DATA_REG_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[15] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_97),
        .Q(\TX_DATA_REG_reg_n_0_[15] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[16] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_96),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[16] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[17] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_95),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[17] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[18] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_94),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[19] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_93),
        .Q(\TX_DATA_REG_reg_n_0_[19] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[1] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(\TX_DATA_REG[1]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[20] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_92),
        .Q(\TX_DATA_REG_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[21] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_91),
        .Q(\TX_DATA_REG_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[22] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_90),
        .Q(\TX_DATA_REG_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[23] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_89),
        .Q(\TX_DATA_REG_reg_n_0_[23] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[24] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_88),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[24] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[25] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_87),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[25] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[26] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_86),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[27] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_85),
        .Q(\TX_DATA_REG_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[28] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_84),
        .Q(\TX_DATA_REG_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[29] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_83),
        .Q(\TX_DATA_REG_reg_n_0_[29] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[2] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_ACK_CNT_n_10),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[30] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_82),
        .Q(\TX_DATA_REG_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[31] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_81),
        .Q(\TX_DATA_REG_reg_n_0_[31] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[32] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_80),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[32] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[33] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_79),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[33] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[34] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_78),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[35] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_77),
        .Q(\TX_DATA_REG_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[36] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_76),
        .Q(\TX_DATA_REG_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[37] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_75),
        .Q(\TX_DATA_REG_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[38] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_74),
        .Q(\TX_DATA_REG_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[39] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_73),
        .Q(\TX_DATA_REG_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[3] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_9),
        .Q(\TX_DATA_REG_reg_n_0_[3] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[40] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_72),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[40] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[41] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_71),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[41] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[42] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_70),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[42] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[43] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_69),
        .Q(\TX_DATA_REG_reg_n_0_[43] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[44] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_68),
        .Q(\TX_DATA_REG_reg_n_0_[44] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[45] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_67),
        .Q(\TX_DATA_REG_reg_n_0_[45] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[46] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_66),
        .Q(\TX_DATA_REG_reg_n_0_[46] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[47] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_65),
        .Q(\TX_DATA_REG_reg_n_0_[47] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[48] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_64),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[48] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[49] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_63),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[49] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[4] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_8),
        .Q(\TX_DATA_REG_reg_n_0_[4] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[50] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_62),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[50] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[51] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_61),
        .Q(\TX_DATA_REG_reg_n_0_[51] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[52] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_60),
        .Q(\TX_DATA_REG_reg_n_0_[52] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[53] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_59),
        .Q(\TX_DATA_REG_reg_n_0_[53] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[54] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_58),
        .Q(\TX_DATA_REG_reg_n_0_[54] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[55] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_57),
        .Q(\TX_DATA_REG_reg_n_0_[55] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[56] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_56),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[56] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[57] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_55),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[57] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[58] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_ACK_CNT_n_4),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[58] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[59] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_3),
        .Q(\TX_DATA_REG_reg_n_0_[59] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[5] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_7),
        .Q(\TX_DATA_REG_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[60] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_54),
        .Q(\TX_DATA_REG_reg_n_0_[60] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[61] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_2),
        .Q(\TX_DATA_REG_reg_n_0_[61] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[62] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_53),
        .Q(\TX_DATA_REG_reg_n_0_[62] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[63] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_1),
        .Q(\TX_DATA_REG_reg_n_0_[63] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[6] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_6),
        .Q(\TX_DATA_REG_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_REG_reg[7] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_5),
        .Q(\TX_DATA_REG_reg_n_0_[7] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[8] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_104),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[8] ));
  FDPE #(
    .INIT(1'b1)) 
    \TX_DATA_REG_reg[9] 
       (.C(clk_i),
        .CE(TX_DATA_REG0),
        .D(U_byte_count_module_n_103),
        .PRE(rst_i),
        .Q(\TX_DATA_REG_reg_n_0_[9] ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[0]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[0]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[0]),
        .Q(\TX_DATA_VALID_DEL11_reg[0]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[1]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[1]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[1]),
        .Q(\TX_DATA_VALID_DEL11_reg[1]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[2]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[2]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[2]),
        .Q(\TX_DATA_VALID_DEL11_reg[2]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[3]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[3]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[3]),
        .Q(\TX_DATA_VALID_DEL11_reg[3]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[4]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[4]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[4]),
        .Q(\TX_DATA_VALID_DEL11_reg[4]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[5]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[5]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[5]),
        .Q(\TX_DATA_VALID_DEL11_reg[5]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[6]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[6]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[6]),
        .Q(\TX_DATA_VALID_DEL11_reg[6]_srl9_activity_blocks_c_7_n_0 ));
  (* srl_bus_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/TX_DATA_VALID_DEL11_reg[7]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \TX_DATA_VALID_DEL11_reg[7]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(TX_DATA_VALID_DEL2[7]),
        .Q(\TX_DATA_VALID_DEL11_reg[7]_srl9_activity_blocks_c_7_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[0]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[0]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[0]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[1]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[1]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[1]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[2]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[2]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[2]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[3]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[3]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[3]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[4]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[4]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[4]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[5]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[5]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[5]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[6]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[6]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[6]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL12_reg[7]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\TX_DATA_VALID_DEL11_reg[7]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\TX_DATA_VALID_DEL12_reg[7]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__7_n_0),
        .Q(TX_DATA_VALID_DEL13__0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__6_n_0),
        .Q(TX_DATA_VALID_DEL13__0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__5_n_0),
        .Q(TX_DATA_VALID_DEL13__0[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__4_n_0),
        .Q(TX_DATA_VALID_DEL13__0[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__3_n_0),
        .Q(TX_DATA_VALID_DEL13__0[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__2_n_0),
        .Q(TX_DATA_VALID_DEL13__0[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__1_n_0),
        .Q(TX_DATA_VALID_DEL13__0[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL13_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate__0_n_0),
        .Q(TX_DATA_VALID_DEL13));
  LUT6 #(
    .INIT(64'hAF0CA300FFFFFFFF)) 
    \TX_DATA_VALID_DEL14[0]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(append_end_frame),
        .I2(txstatplus_int0_out[1]),
        .I3(TX_DATA_VALID_DEL13__0[0]),
        .I4(OVERFLOW_VALID__0[0]),
        .I5(\TX_DATA_VALID_DEL14[0]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL14[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF050DFFFFFFFF)) 
    \TX_DATA_VALID_DEL14[0]_i_2 
       (.I0(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I1(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .I2(TX_DATA_VALID_DEL13__0[0]),
        .I3(fcs_enabled_int),
        .I4(TX_DATA_VALID_DEL13),
        .I5(txstatplus_int0_out[1]),
        .O(\TX_DATA_VALID_DEL14[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAF0CA300FFFFFFFF)) 
    \TX_DATA_VALID_DEL14[1]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(append_end_frame),
        .I2(txstatplus_int0_out[1]),
        .I3(TX_DATA_VALID_DEL13__0[1]),
        .I4(OVERFLOW_VALID__0[1]),
        .I5(\TX_DATA_VALID_DEL14[1]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL14[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF050DFFFFFFFF)) 
    \TX_DATA_VALID_DEL14[1]_i_2 
       (.I0(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I1(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .I2(TX_DATA_VALID_DEL13__0[1]),
        .I3(fcs_enabled_int),
        .I4(TX_DATA_VALID_DEL13),
        .I5(txstatplus_int0_out[1]),
        .O(\TX_DATA_VALID_DEL14[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAF0CA300FFFFFFFF)) 
    \TX_DATA_VALID_DEL14[2]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(append_end_frame),
        .I2(txstatplus_int0_out[1]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .I4(OVERFLOW_VALID__0[2]),
        .I5(\TX_DATA_VALID_DEL14[2]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL14[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0455FFFFFFFF)) 
    \TX_DATA_VALID_DEL14[2]_i_2 
       (.I0(TX_DATA_VALID_DEL13__0[2]),
        .I1(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .I2(fcs_enabled_int),
        .I3(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I4(TX_DATA_VALID_DEL13),
        .I5(txstatplus_int0_out[1]),
        .O(\TX_DATA_VALID_DEL14[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFF0FC50505050)) 
    \TX_DATA_VALID_DEL14[3]_i_1 
       (.I0(\TX_DATA_DEL14[58]_i_6_n_0 ),
        .I1(fcs_enabled_int),
        .I2(TX_DATA_VALID_DEL13__0[3]),
        .I3(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .I4(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14[58]_i_5_n_0 ),
        .O(\TX_DATA_VALID_DEL14[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hCCC0FF3055005500)) 
    \TX_DATA_VALID_DEL14[4]_i_1 
       (.I0(\TX_DATA_DEL14[58]_i_6_n_0 ),
        .I1(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .I2(fcs_enabled_int),
        .I3(TX_DATA_VALID_DEL13__0[4]),
        .I4(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14[58]_i_5_n_0 ),
        .O(\TX_DATA_VALID_DEL14[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair425" *) 
  LUT5 #(
    .INIT(32'hA300FFFF)) 
    \TX_DATA_VALID_DEL14[5]_i_1 
       (.I0(TX_DATA_VALID_DEL13),
        .I1(append_end_frame),
        .I2(txstatplus_int0_out[1]),
        .I3(TX_DATA_VALID_DEL13__0[5]),
        .I4(\TX_DATA_VALID_DEL14[5]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL14[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5D7F557FDDDDDDFF)) 
    \TX_DATA_VALID_DEL14[5]_i_2 
       (.I0(\TX_DATA_DEL14[58]_i_5_n_0 ),
        .I1(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I2(\TX_DATA_VALID_DEL14[7]_i_2_n_0 ),
        .I3(TX_DATA_VALID_DEL13__0[5]),
        .I4(fcs_enabled_int),
        .I5(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DEL14[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0C00FF3055005500)) 
    \TX_DATA_VALID_DEL14[6]_i_1 
       (.I0(\TX_DATA_DEL14[58]_i_6_n_0 ),
        .I1(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ),
        .I2(fcs_enabled_int),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .I4(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I5(\TX_DATA_DEL14[58]_i_5_n_0 ),
        .O(\TX_DATA_VALID_DEL14[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBBFBFFFBFFFFFFFA)) 
    \TX_DATA_VALID_DEL14[6]_i_2 
       (.I0(\TX_DATA_VALID_DEL14[6]_i_3_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[2]),
        .I2(TX_DATA_VALID_DEL13__0[6]),
        .I3(TX_DATA_VALID_DEL13__0[5]),
        .I4(TX_DATA_VALID_DEL13__0[4]),
        .I5(TX_DATA_VALID_DEL13__0[3]),
        .O(\TX_DATA_VALID_DEL14[6]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair441" *) 
  LUT3 #(
    .INIT(8'h7E)) 
    \TX_DATA_VALID_DEL14[6]_i_3 
       (.I0(TX_DATA_VALID_DEL13__0[0]),
        .I1(TX_DATA_VALID_DEL13__0[1]),
        .I2(TX_DATA_VALID_DEL13__0[2]),
        .O(\TX_DATA_VALID_DEL14[6]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair430" *) 
  LUT5 #(
    .INIT(32'hCE00CECC)) 
    \TX_DATA_VALID_DEL14[7]_i_1 
       (.I0(\TX_DATA_VALID_DEL14[7]_i_2_n_0 ),
        .I1(TX_DATA_VALID_DEL13),
        .I2(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ),
        .I3(txstatplus_int0_out[1]),
        .I4(append_end_frame),
        .O(\TX_DATA_VALID_DEL14[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair423" *) 
  LUT5 #(
    .INIT(32'h808A0000)) 
    \TX_DATA_VALID_DEL14[7]_i_2 
       (.I0(\TX_DATA_DEL14[50]_i_5_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[4]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .I4(fcs_enabled_int),
        .O(\TX_DATA_VALID_DEL14[7]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair441" *) 
  LUT4 #(
    .INIT(16'h0051)) 
    \TX_DATA_VALID_DEL14[7]_i_3 
       (.I0(\TX_DATA_VALID_DEL14[7]_i_4_n_0 ),
        .I1(TX_DATA_VALID_DEL13__0[1]),
        .I2(TX_DATA_VALID_DEL13__0[0]),
        .I3(TX_DATA_VALID_DEL13__0[2]),
        .O(\TX_DATA_VALID_DEL14[7]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair422" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \TX_DATA_VALID_DEL14[7]_i_4 
       (.I0(TX_DATA_VALID_DEL13__0[3]),
        .I1(TX_DATA_VALID_DEL13__0[4]),
        .I2(TX_DATA_VALID_DEL13__0[5]),
        .I3(TX_DATA_VALID_DEL13__0[6]),
        .O(\TX_DATA_VALID_DEL14[7]_i_4_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[0]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[1]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[2]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[3]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[4]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[5]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[6]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL14_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_DEL14[7]_i_1_n_0 ),
        .Q(TX_DATA_VALID_DEL14[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[0]),
        .Q(TX_DATA_VALID_DEL15[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[1]),
        .Q(TX_DATA_VALID_DEL15[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[2]),
        .Q(TX_DATA_VALID_DEL15[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[3]),
        .Q(TX_DATA_VALID_DEL15[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[4]),
        .Q(TX_DATA_VALID_DEL15[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[5]),
        .Q(TX_DATA_VALID_DEL15[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[6]),
        .Q(TX_DATA_VALID_DEL15[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL15_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL14[7]),
        .Q(TX_DATA_VALID_DEL15[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[0] ),
        .Q(TX_DATA_VALID_DEL1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[1] ),
        .Q(TX_DATA_VALID_DEL1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[2] ),
        .Q(TX_DATA_VALID_DEL1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[3] ),
        .Q(TX_DATA_VALID_DEL1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[4] ),
        .Q(TX_DATA_VALID_DEL1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[5] ),
        .Q(TX_DATA_VALID_DEL1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[6] ),
        .Q(TX_DATA_VALID_DEL1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\TX_DATA_VALID_REG_reg_n_0_[7] ),
        .Q(TX_DATA_VALID_DEL1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[0]),
        .Q(TX_DATA_VALID_DEL2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[1]),
        .Q(TX_DATA_VALID_DEL2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[2]),
        .Q(TX_DATA_VALID_DEL2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[3]),
        .Q(TX_DATA_VALID_DEL2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[4]),
        .Q(TX_DATA_VALID_DEL2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[5]),
        .Q(TX_DATA_VALID_DEL2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[6]),
        .Q(TX_DATA_VALID_DEL2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DEL2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL1[7]),
        .Q(TX_DATA_VALID_DEL2[7]));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[0]),
        .Q(TX_DATA_VALID_DELAY[0]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[10]),
        .Q(TX_DATA_VALID_DELAY[10]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[11]),
        .Q(TX_DATA_VALID_DELAY[11]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[12]),
        .Q(TX_DATA_VALID_DELAY[12]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[13]),
        .Q(TX_DATA_VALID_DELAY[13]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[14]),
        .Q(TX_DATA_VALID_DELAY[14]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[15]),
        .Q(TX_DATA_VALID_DELAY[15]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[16]),
        .Q(TX_DATA_VALID_DELAY[16]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[17]),
        .Q(TX_DATA_VALID_DELAY[17]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[18]),
        .Q(TX_DATA_VALID_DELAY[18]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[19]),
        .Q(TX_DATA_VALID_DELAY[19]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[1]),
        .Q(TX_DATA_VALID_DELAY[1]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[20]),
        .Q(TX_DATA_VALID_DELAY[20]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[21]),
        .Q(TX_DATA_VALID_DELAY[21]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[22]),
        .Q(TX_DATA_VALID_DELAY[22]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[23]),
        .Q(TX_DATA_VALID_DELAY[23]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[24]),
        .Q(TX_DATA_VALID_DELAY[24]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[25]),
        .Q(TX_DATA_VALID_DELAY[25]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[26]),
        .Q(TX_DATA_VALID_DELAY[26]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[27]),
        .Q(TX_DATA_VALID_DELAY[27]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[28]),
        .Q(TX_DATA_VALID_DELAY[28]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[29]),
        .Q(TX_DATA_VALID_DELAY[29]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[2]),
        .Q(TX_DATA_VALID_DELAY[2]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[30]),
        .Q(TX_DATA_VALID_DELAY[30]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[31]),
        .Q(TX_DATA_VALID_DELAY[31]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[32]),
        .Q(TX_DATA_VALID_DELAY[32]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[33]),
        .Q(TX_DATA_VALID_DELAY[33]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[34]),
        .Q(TX_DATA_VALID_DELAY[34]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[35]),
        .Q(TX_DATA_VALID_DELAY[35]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[36]),
        .Q(TX_DATA_VALID_DELAY[36]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[37]),
        .Q(TX_DATA_VALID_DELAY[37]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[38]),
        .Q(TX_DATA_VALID_DELAY[38]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[39]),
        .Q(TX_DATA_VALID_DELAY[39]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[3]),
        .Q(TX_DATA_VALID_DELAY[3]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[40]),
        .Q(TX_DATA_VALID_DELAY[40]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[41]),
        .Q(TX_DATA_VALID_DELAY[41]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[42]),
        .Q(TX_DATA_VALID_DELAY[42]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[43]),
        .Q(TX_DATA_VALID_DELAY[43]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[44]),
        .Q(TX_DATA_VALID_DELAY[44]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[45]),
        .Q(TX_DATA_VALID_DELAY[45]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[46]),
        .Q(TX_DATA_VALID_DELAY[46]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[47]),
        .Q(TX_DATA_VALID_DELAY[47]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[48]),
        .Q(TX_DATA_VALID_DELAY[48]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[49]),
        .Q(TX_DATA_VALID_DELAY[49]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[4]),
        .Q(TX_DATA_VALID_DELAY[4]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[50]),
        .Q(TX_DATA_VALID_DELAY[50]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[51]),
        .Q(TX_DATA_VALID_DELAY[51]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[52]),
        .Q(TX_DATA_VALID_DELAY[52]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[53]),
        .Q(TX_DATA_VALID_DELAY[53]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[54]),
        .Q(TX_DATA_VALID_DELAY[54]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[55]),
        .Q(TX_DATA_VALID_DELAY[55]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[56]),
        .Q(TX_DATA_VALID_DELAY[56]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[57]),
        .Q(TX_DATA_VALID_DELAY[57]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[58]),
        .Q(TX_DATA_VALID_DELAY[58]),
        .S(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[59]),
        .Q(TX_DATA_VALID_DELAY[59]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[5]),
        .Q(TX_DATA_VALID_DELAY[5]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[60]),
        .Q(TX_DATA_VALID_DELAY[60]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[61]),
        .Q(TX_DATA_VALID_DELAY[61]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[62]),
        .Q(TX_DATA_VALID_DELAY[62]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[63]),
        .Q(TX_DATA_VALID_DELAY[63]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[6]),
        .Q(TX_DATA_VALID_DELAY[6]),
        .R(out));
  FDRE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_DELAY_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[7]),
        .Q(TX_DATA_VALID_DELAY[7]),
        .R(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[8]),
        .Q(TX_DATA_VALID_DELAY[8]),
        .S(out));
  FDSE #(
    .INIT(1'b1)) 
    \TX_DATA_VALID_DELAY_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(TX_DATA[9]),
        .Q(TX_DATA_VALID_DELAY[9]),
        .S(out));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_52),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_51),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_50),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_49),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_48),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_47),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_46),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \TX_DATA_VALID_REG_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(U_byte_count_module_n_45),
        .Q(\TX_DATA_VALID_REG_reg_n_0_[7] ));
  FDRE #(
    .INIT(1'b0)) 
    TX_STATS_VALID_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(append_end_frame),
        .Q(TX_STATS_VALID),
        .R(1'b0));
  switch_elements_ack_counter U_ACK_CNT
       (.AR(RESET02_out),
        .D({U_ACK_CNT_n_1,U_ACK_CNT_n_2,U_ACK_CNT_n_3,U_ACK_CNT_n_4,U_ACK_CNT_n_5,U_ACK_CNT_n_6,U_ACK_CNT_n_7,U_ACK_CNT_n_8,U_ACK_CNT_n_9,U_ACK_CNT_n_10}),
        .E(U_ACK_CNT_n_13),
        .\FC_TX_PAUSEDATA_reg[15] ({U_ACK_CNT_n_24,U_ACK_CNT_n_25,U_ACK_CNT_n_26,U_ACK_CNT_n_27,U_ACK_CNT_n_28,U_ACK_CNT_n_29,U_ACK_CNT_n_30,U_ACK_CNT_n_31,U_ACK_CNT_n_32,U_ACK_CNT_n_33,U_ACK_CNT_n_34,U_ACK_CNT_n_35,U_ACK_CNT_n_36,U_ACK_CNT_n_37,U_ACK_CNT_n_38,U_ACK_CNT_n_39}),
        .FRAME_START(FRAME_START),
        .I94(I94),
        .Q(DELAY_ACK),
        .SS(RESET0),
        .\TX_DATA_REG_reg[40] ({shift_pause_data[56],shift_pause_data[15],shift_pause_data[13],shift_pause_data[11:10],shift_pause_data[8:2]}),
        .\TX_DATA_REG_reg[63] (U_byte_count_module_n_105),
        .\TX_DATA_REG_reg[63]_0 ({\TX_DATA_VALID_REG_reg_n_0_[7] ,\TX_DATA_VALID_REG_reg_n_0_[0] }),
        .\TX_DATA_REG_reg[63]_1 ({TX_DATA_VALID_DELAY[63],TX_DATA_VALID_DELAY[61],TX_DATA_VALID_DELAY[59:58],TX_DATA_VALID_DELAY[7:2]}),
        .append_start_pause(append_start_pause),
        .append_start_pause_reg(U_ACK_CNT_n_11),
        .append_start_pause_reg_0(U_ACK_CNT_n_12),
        .apply_pause_delay(apply_pause_delay),
        .apply_pause_delay_reg(apply_pause_delay_reg_0),
        .clk_i(clk_i),
        .out(out),
        .reset_tx_int(reset_tx_int),
        .rst_i(rst_i),
        .start_count_del_reg_0(transmit_pause_frame_reg_n_0),
        .transmit_pause_frame_valid(transmit_pause_frame_valid),
        .tx_ack_reg_0(TX_ACK),
        .tx_ack_reg_1(U_ACK_CNT_n_16),
        .tx_ack_reg_2(U_ACK_CNT_n_17),
        .tx_ack_reg_3(U_ACK_CNT_n_18),
        .tx_ack_reg_4(U_ACK_CNT_n_19),
        .tx_ack_reg_5(U_ACK_CNT_n_20),
        .tx_ack_reg_6(U_ACK_CNT_n_21),
        .tx_ack_reg_7(U_ACK_CNT_n_22));
  switch_elements_CRC32_D64 U_CRC64
       (.\CRC_OUT_reg[24]_0 ({\TX_DATA_REG_reg_n_0_[63] ,\TX_DATA_REG_reg_n_0_[62] ,\TX_DATA_REG_reg_n_0_[61] ,\TX_DATA_REG_reg_n_0_[60] ,\TX_DATA_REG_reg_n_0_[59] ,\TX_DATA_REG_reg_n_0_[58] ,\TX_DATA_REG_reg_n_0_[57] ,\TX_DATA_REG_reg_n_0_[56] ,\TX_DATA_REG_reg_n_0_[55] ,\TX_DATA_REG_reg_n_0_[54] ,\TX_DATA_REG_reg_n_0_[53] ,\TX_DATA_REG_reg_n_0_[52] ,\TX_DATA_REG_reg_n_0_[51] ,\TX_DATA_REG_reg_n_0_[50] ,\TX_DATA_REG_reg_n_0_[49] ,\TX_DATA_REG_reg_n_0_[48] ,\TX_DATA_REG_reg_n_0_[47] ,\TX_DATA_REG_reg_n_0_[46] ,\TX_DATA_REG_reg_n_0_[45] ,\TX_DATA_REG_reg_n_0_[44] ,\TX_DATA_REG_reg_n_0_[43] ,\TX_DATA_REG_reg_n_0_[42] ,\TX_DATA_REG_reg_n_0_[41] ,\TX_DATA_REG_reg_n_0_[40] ,\TX_DATA_REG_reg_n_0_[39] ,\TX_DATA_REG_reg_n_0_[38] ,\TX_DATA_REG_reg_n_0_[37] ,\TX_DATA_REG_reg_n_0_[36] ,\TX_DATA_REG_reg_n_0_[35] ,\TX_DATA_REG_reg_n_0_[34] ,\TX_DATA_REG_reg_n_0_[33] ,\TX_DATA_REG_reg_n_0_[32] ,\TX_DATA_REG_reg_n_0_[31] ,\TX_DATA_REG_reg_n_0_[30] ,\TX_DATA_REG_reg_n_0_[29] ,\TX_DATA_REG_reg_n_0_[28] ,\TX_DATA_REG_reg_n_0_[27] ,\TX_DATA_REG_reg_n_0_[26] ,\TX_DATA_REG_reg_n_0_[25] ,\TX_DATA_REG_reg_n_0_[24] ,\TX_DATA_REG_reg_n_0_[23] ,\TX_DATA_REG_reg_n_0_[22] ,\TX_DATA_REG_reg_n_0_[21] ,\TX_DATA_REG_reg_n_0_[20] ,\TX_DATA_REG_reg_n_0_[19] ,\TX_DATA_REG_reg_n_0_[18] ,\TX_DATA_REG_reg_n_0_[17] ,\TX_DATA_REG_reg_n_0_[16] ,\TX_DATA_REG_reg_n_0_[15] ,\TX_DATA_REG_reg_n_0_[14] ,\TX_DATA_REG_reg_n_0_[13] ,\TX_DATA_REG_reg_n_0_[12] ,\TX_DATA_REG_reg_n_0_[11] ,\TX_DATA_REG_reg_n_0_[10] ,\TX_DATA_REG_reg_n_0_[9] ,\TX_DATA_REG_reg_n_0_[8] ,\TX_DATA_REG_reg_n_0_[7] ,\TX_DATA_REG_reg_n_0_[6] ,\TX_DATA_REG_reg_n_0_[5] ,\TX_DATA_REG_reg_n_0_[4] ,\TX_DATA_REG_reg_n_0_[3] ,\TX_DATA_REG_reg_n_0_[2] ,\TX_DATA_REG_reg_n_0_[1] ,\TX_DATA_REG_reg_n_0_[0] }),
        .Q(CRC_32_64),
        .SS(RESET0),
        .clk_i(clk_i),
        .frame_start_del(frame_start_del),
        .transmit_pause_frame_valid(transmit_pause_frame_valid));
  switch_elements_CRC32_D8 U_CRC8
       (.\CRC_OUT_reg[31]_0 (CRC_32_64),
        .D({U_CRC8_n_0,U_CRC8_n_1,U_CRC8_n_2,U_CRC8_n_3,U_CRC8_n_4,U_CRC8_n_5,U_CRC8_n_6,U_CRC8_n_7,U_CRC8_n_8,U_CRC8_n_9,U_CRC8_n_10,U_CRC8_n_11,U_CRC8_n_12,U_CRC8_n_13,U_CRC8_n_14,U_CRC8_n_15,U_CRC8_n_16,U_CRC8_n_17,U_CRC8_n_18,U_CRC8_n_19,U_CRC8_n_20,U_CRC8_n_21,U_CRC8_n_22,U_CRC8_n_23}),
        .E(U_CRC8_n_24),
        .\OVERFLOW_DATA_reg[19] (\OVERFLOW_DATA[23]_i_2_n_0 ),
        .\OVERFLOW_DATA_reg[2] (\OVERFLOW_DATA[31]_i_2_n_0 ),
        .\OVERFLOW_DATA_reg[2]_0 (\OVERFLOW_DATA[17]_i_2_n_0 ),
        .\OVERFLOW_DATA_reg[8] (\OVERFLOW_DATA[8]_i_2_n_0 ),
        .Q(tx_data_int),
        .TX_DATA_DEL13(TX_DATA_DEL13),
        .\TX_DATA_DEL14[57]_i_2_0 (\TX_DATA_DEL14[57]_i_8_n_0 ),
        .\TX_DATA_DEL14[57]_i_2_1 (\TX_DATA_DEL14[57]_i_7_n_0 ),
        .\TX_DATA_DEL14[57]_i_2_2 (\TX_DATA_VALID_DEL14[6]_i_3_n_0 ),
        .\TX_DATA_DEL14[63]_i_2_0 (\TX_DATA_DEL14[50]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[0] (\TX_DATA_DEL14[15]_i_2_n_0 ),
        .\TX_DATA_DEL14_reg[18] (\TX_DATA_DEL14[23]_i_2_n_0 ),
        .\TX_DATA_DEL14_reg[18]_0 (\TX_DATA_DEL14[18]_i_4_n_0 ),
        .\TX_DATA_DEL14_reg[21] (\TX_DATA_DEL14[63]_i_7_n_0 ),
        .\TX_DATA_DEL14_reg[25] (\TX_DATA_DEL14[25]_i_4_n_0 ),
        .\TX_DATA_DEL14_reg[26] (\TX_DATA_DEL14[39]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[32] (\TX_DATA_DEL14[63]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[32]_0 (\TX_DATA_DEL14[63]_i_4_n_0 ),
        .\TX_DATA_DEL14_reg[33] (\TX_DATA_DEL14[33]_i_6_n_0 ),
        .\TX_DATA_DEL14_reg[33]_0 (\TX_DATA_DEL14[33]_i_4_n_0 ),
        .\TX_DATA_DEL14_reg[38] ({\OVERFLOW_DATA_reg_n_0_[39] ,\OVERFLOW_DATA_reg_n_0_[33] ,\OVERFLOW_DATA_reg_n_0_[31] ,\OVERFLOW_DATA_reg_n_0_[23] ,\OVERFLOW_DATA_reg_n_0_[22] ,\OVERFLOW_DATA_reg_n_0_[21] ,\OVERFLOW_DATA_reg_n_0_[20] ,\OVERFLOW_DATA_reg_n_0_[19] ,\OVERFLOW_DATA_reg_n_0_[17] ,\OVERFLOW_DATA_reg_n_0_[16] ,\OVERFLOW_DATA_reg_n_0_[15] ,\OVERFLOW_DATA_reg_n_0_[14] ,\OVERFLOW_DATA_reg_n_0_[13] ,\OVERFLOW_DATA_reg_n_0_[12] ,\OVERFLOW_DATA_reg_n_0_[11] ,\OVERFLOW_DATA_reg_n_0_[10] ,\OVERFLOW_DATA_reg_n_0_[9] ,\OVERFLOW_DATA_reg_n_0_[8] ,\OVERFLOW_DATA_reg_n_0_[7] ,\OVERFLOW_DATA_reg_n_0_[6] ,\OVERFLOW_DATA_reg_n_0_[5] ,\OVERFLOW_DATA_reg_n_0_[4] ,\OVERFLOW_DATA_reg_n_0_[3] ,\OVERFLOW_DATA_reg_n_0_[2] ,\OVERFLOW_DATA_reg_n_0_[1] ,\OVERFLOW_DATA_reg_n_0_[0] }),
        .\TX_DATA_DEL14_reg[39] (\TX_DATA_DEL14[39]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[41] (\TX_DATA_DEL14[41]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[47] (\TX_DATA_DEL14[47]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[48] (\TX_DATA_DEL14[48]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[48]_0 (\TX_DATA_DEL14[48]_i_6_n_0 ),
        .\TX_DATA_DEL14_reg[49] (\TX_DATA_DEL14[49]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[49]_0 (\TX_DATA_DEL14[49]_i_6_n_0 ),
        .\TX_DATA_DEL14_reg[50] (\TX_DATA_DEL14[50]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[51] (\TX_DATA_DEL14[51]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[52] (\TX_DATA_DEL14[52]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[53] (\TX_DATA_DEL14[53]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[54] (\TX_DATA_DEL14[54]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[54]_0 (\TX_DATA_DEL14[54]_i_6_n_0 ),
        .\TX_DATA_DEL14_reg[55] (\TX_DATA_DEL14[55]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[57] (\TX_DATA_DEL14[57]_i_6_n_0 ),
        .\TX_DATA_DEL14_reg[58] (\TX_DATA_DEL14[58]_i_3_n_0 ),
        .\TX_DATA_DEL14_reg[58]_0 (\TX_DATA_DEL14[58]_i_5_n_0 ),
        .\TX_DATA_DEL14_reg[58]_1 (\TX_DATA_DEL14[58]_i_6_n_0 ),
        .TX_DATA_VALID_DEL13(TX_DATA_VALID_DEL13),
        .TX_DATA_VALID_DEL13__0({TX_DATA_VALID_DEL13__0[6:4],TX_DATA_VALID_DEL13__0[2:0]}),
        .\TX_DATA_VALID_DEL13_reg[7] ({U_CRC8_n_25,U_CRC8_n_26,U_CRC8_n_27,U_CRC8_n_28,U_CRC8_n_29,U_CRC8_n_30,U_CRC8_n_31,U_CRC8_n_32,U_CRC8_n_33,U_CRC8_n_34,U_CRC8_n_35,U_CRC8_n_36,U_CRC8_n_37,U_CRC8_n_38,U_CRC8_n_39,U_CRC8_n_40,U_CRC8_n_41,U_CRC8_n_42,U_CRC8_n_43,U_CRC8_n_44,U_CRC8_n_45,U_CRC8_n_46,U_CRC8_n_47,U_CRC8_n_48,U_CRC8_n_49,U_CRC8_n_50,U_CRC8_n_51,U_CRC8_n_52,U_CRC8_n_53,U_CRC8_n_54,U_CRC8_n_55,U_CRC8_n_56,U_CRC8_n_57,U_CRC8_n_58,U_CRC8_n_59,U_CRC8_n_60,U_CRC8_n_61,U_CRC8_n_62,U_CRC8_n_63,U_CRC8_n_64,U_CRC8_n_65,U_CRC8_n_66,U_CRC8_n_67,U_CRC8_n_68,U_CRC8_n_69,U_CRC8_n_70,U_CRC8_n_71,U_CRC8_n_72,U_CRC8_n_73,U_CRC8_n_74,U_CRC8_n_75,U_CRC8_n_76,U_CRC8_n_77,U_CRC8_n_78,U_CRC8_n_79,U_CRC8_n_80,U_CRC8_n_81,U_CRC8_n_82,U_CRC8_n_83,U_CRC8_n_84,U_CRC8_n_85,U_CRC8_n_86,U_CRC8_n_87,U_CRC8_n_88}),
        .append_end_frame(append_end_frame),
        .clk_i(clk_i),
        .fcs_enabled_int(fcs_enabled_int),
        .load_CRC8(load_CRC8),
        .rst_i(rst_i),
        .start_CRC8(start_CRC8),
        .txstatplus_int(txstatplus_int),
        .txstatplus_int0_out(txstatplus_int0_out[1]));
  switch_elements_byte_count_module U_byte_count_module
       (.AR(RESET02_out),
        .\BYTE_COUNTER_reg[3]_0 (U_byte_count_module_n_105),
        .\BYTE_COUNTER_reg[3]_1 (TX_DATA_REG0),
        .D(p_0_in__2[15:2]),
        .E(length_register0),
        .FRAME_START(FRAME_START),
        .FRAME_START_reg(FRAME_START_i_3_n_0),
        .Q(BYTE_COUNTER),
        .TX_ACK(TX_ACK),
        .\TX_DATA_REG_reg[0] (\TX_DATA_REG[63]_i_4_n_0 ),
        .\TX_DATA_REG_reg[10] (U_ACK_CNT_n_17),
        .\TX_DATA_REG_reg[11] (U_ACK_CNT_n_19),
        .\TX_DATA_REG_reg[12] (\TX_DATA_REG[12]_i_2_n_0 ),
        .\TX_DATA_REG_reg[13] (U_ACK_CNT_n_20),
        .\TX_DATA_REG_reg[14] (\TX_DATA_REG[14]_i_2_n_0 ),
        .\TX_DATA_REG_reg[15] ({U_byte_count_module_n_28,U_byte_count_module_n_29,U_byte_count_module_n_30,U_byte_count_module_n_31,U_byte_count_module_n_32,U_byte_count_module_n_33,U_byte_count_module_n_34,U_byte_count_module_n_35,U_byte_count_module_n_36,U_byte_count_module_n_37,U_byte_count_module_n_38,U_byte_count_module_n_39,U_byte_count_module_n_40,U_byte_count_module_n_41,U_byte_count_module_n_42,U_byte_count_module_n_43}),
        .\TX_DATA_REG_reg[15]_0 (U_ACK_CNT_n_21),
        .\TX_DATA_REG_reg[16] (U_ACK_CNT_n_12),
        .\TX_DATA_REG_reg[19] (U_ACK_CNT_n_22),
        .\TX_DATA_REG_reg[20] (\TX_DATA_REG[60]_i_2_n_0 ),
        .\TX_DATA_REG_reg[21] (U_ACK_CNT_n_11),
        .\TX_DATA_REG_reg[33] (\TX_DATA_REG[56]_i_2_n_0 ),
        .\TX_DATA_REG_reg[40] (U_ACK_CNT_n_18),
        .\TX_DATA_REG_reg[62] ({\TX_DATA_VALID_REG_reg_n_0_[7] ,\TX_DATA_VALID_REG_reg_n_0_[6] ,\TX_DATA_VALID_REG_reg_n_0_[5] ,\TX_DATA_VALID_REG_reg_n_0_[4] ,\TX_DATA_VALID_REG_reg_n_0_[3] ,\TX_DATA_VALID_REG_reg_n_0_[2] ,\TX_DATA_VALID_REG_reg_n_0_[1] ,\TX_DATA_VALID_REG_reg_n_0_[0] }),
        .\TX_DATA_REG_reg[62]_0 ({TX_DATA_VALID_DELAY[62],TX_DATA_VALID_DELAY[60],TX_DATA_VALID_DELAY[57:8]}),
        .\TX_DATA_REG_reg[8] (U_ACK_CNT_n_16),
        .\TX_DATA_REG_reg[9] (\TX_DATA_REG[9]_i_2_n_0 ),
        .\TX_DATA_VALID_DELAY_reg[62] ({U_byte_count_module_n_53,U_byte_count_module_n_54,U_byte_count_module_n_55,U_byte_count_module_n_56,U_byte_count_module_n_57,U_byte_count_module_n_58,U_byte_count_module_n_59,U_byte_count_module_n_60,U_byte_count_module_n_61,U_byte_count_module_n_62,U_byte_count_module_n_63,U_byte_count_module_n_64,U_byte_count_module_n_65,U_byte_count_module_n_66,U_byte_count_module_n_67,U_byte_count_module_n_68,U_byte_count_module_n_69,U_byte_count_module_n_70,U_byte_count_module_n_71,U_byte_count_module_n_72,U_byte_count_module_n_73,U_byte_count_module_n_74,U_byte_count_module_n_75,U_byte_count_module_n_76,U_byte_count_module_n_77,U_byte_count_module_n_78,U_byte_count_module_n_79,U_byte_count_module_n_80,U_byte_count_module_n_81,U_byte_count_module_n_82,U_byte_count_module_n_83,U_byte_count_module_n_84,U_byte_count_module_n_85,U_byte_count_module_n_86,U_byte_count_module_n_87,U_byte_count_module_n_88,U_byte_count_module_n_89,U_byte_count_module_n_90,U_byte_count_module_n_91,U_byte_count_module_n_92,U_byte_count_module_n_93,U_byte_count_module_n_94,U_byte_count_module_n_95,U_byte_count_module_n_96,U_byte_count_module_n_97,U_byte_count_module_n_98,U_byte_count_module_n_99,U_byte_count_module_n_100,U_byte_count_module_n_101,U_byte_count_module_n_102,U_byte_count_module_n_103,U_byte_count_module_n_104}),
        .\TX_DATA_VALID_REG_reg[4] ({shift_pause_valid_del[4],shift_pause_valid_del[0]}),
        .\TX_DATA_VALID_REG_reg[7] (\TX_DATA_VALID_REG_reg[7]_0 ),
        .clk_i(clk_i),
        .\enable_i[6] ({U_byte_count_module_n_45,U_byte_count_module_n_46,U_byte_count_module_n_47,U_byte_count_module_n_48,U_byte_count_module_n_49,U_byte_count_module_n_50,U_byte_count_module_n_51,U_byte_count_module_n_52}),
        .\final_byte_count_reg[10] (\final_byte_count[10]_i_2_n_0 ),
        .\final_byte_count_reg[11] (\final_byte_count[12]_i_2_n_0 ),
        .\final_byte_count_reg[13] (\final_byte_count[13]_i_2_n_0 ),
        .\final_byte_count_reg[14] (\final_byte_count[15]_i_3_n_0 ),
        .\final_byte_count_reg[15] (byte_count_reg),
        .\final_byte_count_reg[15]_0 ({final_byte_count_reg__0,final_byte_count_reg}),
        .\final_byte_count_reg[3] (\final_byte_count[3]_i_2_n_0 ),
        .\final_byte_count_reg[4] (\final_byte_count[4]_i_2_n_0 ),
        .\final_byte_count_reg[5] (\final_byte_count[5]_i_3_n_0 ),
        .\final_byte_count_reg[6] (\final_byte_count[7]_i_2_n_0 ),
        .\final_byte_count_reg[8] (\final_byte_count[8]_i_2_n_0 ),
        .\final_byte_count_reg[9] (\final_byte_count[9]_i_2_n_0 ),
        .frame_start_del(frame_start_del),
        .\length_register_reg[15] ({\TX_DATA_REG_reg_n_0_[47] ,\TX_DATA_REG_reg_n_0_[46] ,\TX_DATA_REG_reg_n_0_[45] ,\TX_DATA_REG_reg_n_0_[44] ,\TX_DATA_REG_reg_n_0_[43] ,\TX_DATA_REG_reg_n_0_[42] ,\TX_DATA_REG_reg_n_0_[41] ,\TX_DATA_REG_reg_n_0_[40] ,\TX_DATA_REG_reg_n_0_[39] ,\TX_DATA_REG_reg_n_0_[38] ,\TX_DATA_REG_reg_n_0_[37] ,\TX_DATA_REG_reg_n_0_[36] ,\TX_DATA_REG_reg_n_0_[35] ,\TX_DATA_REG_reg_n_0_[34] ,\TX_DATA_REG_reg_n_0_[33] ,\TX_DATA_REG_reg_n_0_[32] ,\TX_DATA_REG_reg_n_0_[15] ,\TX_DATA_REG_reg_n_0_[14] ,\TX_DATA_REG_reg_n_0_[13] ,\TX_DATA_REG_reg_n_0_[12] ,\TX_DATA_REG_reg_n_0_[11] ,\TX_DATA_REG_reg_n_0_[10] ,\TX_DATA_REG_reg_n_0_[9] ,\TX_DATA_REG_reg_n_0_[8] ,\TX_DATA_REG_reg_n_0_[7] ,\TX_DATA_REG_reg_n_0_[6] ,\TX_DATA_REG_reg_n_0_[5] ,\TX_DATA_REG_reg_n_0_[4] ,\TX_DATA_REG_reg_n_0_[3] ,\TX_DATA_REG_reg_n_0_[2] ,\TX_DATA_REG_reg_n_0_[1] ,\TX_DATA_REG_reg_n_0_[0] }),
        .load_CRC8(load_CRC8),
        .out(out),
        .transmit_pause_frame_del(transmit_pause_frame_del),
        .transmit_pause_frame_valid(transmit_pause_frame_valid),
        .tx_ack_reg(U_byte_count_module_n_107),
        .vlan_enabled_int(vlan_enabled_int));
  (* SOFT_HLUTNM = "soft_lutpair492" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate
       (.I0(\append_reg_reg[9]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate_n_0));
  (* SOFT_HLUTNM = "soft_lutpair493" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__0
       (.I0(\TX_DATA_VALID_DEL12_reg[7]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair494" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__1
       (.I0(\TX_DATA_VALID_DEL12_reg[6]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair503" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__10
       (.I0(\TX_DATA_DEL12_reg[61]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair504" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__11
       (.I0(\TX_DATA_DEL12_reg[60]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__11_n_0));
  (* SOFT_HLUTNM = "soft_lutpair505" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__12
       (.I0(\TX_DATA_DEL12_reg[59]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair507" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__13
       (.I0(\TX_DATA_DEL12_reg[58]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__13_n_0));
  (* SOFT_HLUTNM = "soft_lutpair508" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__14
       (.I0(\TX_DATA_DEL12_reg[57]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__14_n_0));
  (* SOFT_HLUTNM = "soft_lutpair509" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__15
       (.I0(\TX_DATA_DEL12_reg[56]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair510" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__16
       (.I0(\TX_DATA_DEL12_reg[55]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair511" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__17
       (.I0(\TX_DATA_DEL12_reg[54]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair512" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__18
       (.I0(\TX_DATA_DEL12_reg[53]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair513" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__19
       (.I0(\TX_DATA_DEL12_reg[52]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__19_n_0));
  (* SOFT_HLUTNM = "soft_lutpair495" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__2
       (.I0(\TX_DATA_VALID_DEL12_reg[5]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair514" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__20
       (.I0(\TX_DATA_DEL12_reg[51]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__20_n_0));
  (* SOFT_HLUTNM = "soft_lutpair517" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__21
       (.I0(\TX_DATA_DEL12_reg[50]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__21_n_0));
  (* SOFT_HLUTNM = "soft_lutpair518" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__22
       (.I0(\TX_DATA_DEL12_reg[49]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__22_n_0));
  (* SOFT_HLUTNM = "soft_lutpair519" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__23
       (.I0(\TX_DATA_DEL12_reg[48]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__23_n_0));
  (* SOFT_HLUTNM = "soft_lutpair520" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__24
       (.I0(\TX_DATA_DEL12_reg[47]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__24_n_0));
  (* SOFT_HLUTNM = "soft_lutpair521" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__25
       (.I0(\TX_DATA_DEL12_reg[46]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__25_n_0));
  (* SOFT_HLUTNM = "soft_lutpair522" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__26
       (.I0(\TX_DATA_DEL12_reg[45]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__26_n_0));
  (* SOFT_HLUTNM = "soft_lutpair523" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__27
       (.I0(\TX_DATA_DEL12_reg[44]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__27_n_0));
  (* SOFT_HLUTNM = "soft_lutpair524" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__28
       (.I0(\TX_DATA_DEL12_reg[43]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__28_n_0));
  (* SOFT_HLUTNM = "soft_lutpair525" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__29
       (.I0(\TX_DATA_DEL12_reg[42]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__29_n_0));
  (* SOFT_HLUTNM = "soft_lutpair496" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__3
       (.I0(\TX_DATA_VALID_DEL12_reg[4]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__3_n_0));
  (* SOFT_HLUTNM = "soft_lutpair526" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__30
       (.I0(\TX_DATA_DEL12_reg[41]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__30_n_0));
  (* SOFT_HLUTNM = "soft_lutpair526" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__31
       (.I0(\TX_DATA_DEL12_reg[40]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__31_n_0));
  (* SOFT_HLUTNM = "soft_lutpair527" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__32
       (.I0(\TX_DATA_DEL12_reg[39]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__32_n_0));
  (* SOFT_HLUTNM = "soft_lutpair527" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__33
       (.I0(\TX_DATA_DEL12_reg[38]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__33_n_0));
  (* SOFT_HLUTNM = "soft_lutpair528" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__34
       (.I0(\TX_DATA_DEL12_reg[37]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__34_n_0));
  (* SOFT_HLUTNM = "soft_lutpair528" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__35
       (.I0(\TX_DATA_DEL12_reg[36]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__35_n_0));
  (* SOFT_HLUTNM = "soft_lutpair536" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__36
       (.I0(\TX_DATA_DEL12_reg[35]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__36_n_0));
  (* SOFT_HLUTNM = "soft_lutpair536" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__37
       (.I0(\TX_DATA_DEL12_reg[34]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__37_n_0));
  (* SOFT_HLUTNM = "soft_lutpair537" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__38
       (.I0(\TX_DATA_DEL12_reg[33]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__38_n_0));
  (* SOFT_HLUTNM = "soft_lutpair525" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__39
       (.I0(\TX_DATA_DEL12_reg[32]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__39_n_0));
  (* SOFT_HLUTNM = "soft_lutpair497" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__4
       (.I0(\TX_DATA_VALID_DEL12_reg[3]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__4_n_0));
  (* SOFT_HLUTNM = "soft_lutpair524" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__40
       (.I0(\TX_DATA_DEL12_reg[31]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__40_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__41
       (.I0(\TX_DATA_DEL12_reg[30]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__41_n_0));
  (* SOFT_HLUTNM = "soft_lutpair512" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__42
       (.I0(\TX_DATA_DEL12_reg[29]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__42_n_0));
  (* SOFT_HLUTNM = "soft_lutpair504" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__43
       (.I0(\TX_DATA_DEL12_reg[28]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__43_n_0));
  (* SOFT_HLUTNM = "soft_lutpair503" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__44
       (.I0(\TX_DATA_DEL12_reg[27]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__44_n_0));
  (* SOFT_HLUTNM = "soft_lutpair502" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__45
       (.I0(\TX_DATA_DEL12_reg[26]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__45_n_0));
  (* SOFT_HLUTNM = "soft_lutpair518" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__46
       (.I0(\TX_DATA_DEL12_reg[25]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__46_n_0));
  (* SOFT_HLUTNM = "soft_lutpair537" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__47
       (.I0(\TX_DATA_DEL12_reg[24]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__47_n_0));
  (* SOFT_HLUTNM = "soft_lutpair499" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__48
       (.I0(\TX_DATA_DEL12_reg[23]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__48_n_0));
  (* SOFT_HLUTNM = "soft_lutpair514" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__49
       (.I0(\TX_DATA_DEL12_reg[22]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__49_n_0));
  (* SOFT_HLUTNM = "soft_lutpair498" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__5
       (.I0(\TX_DATA_VALID_DEL12_reg[2]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair513" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__50
       (.I0(\TX_DATA_DEL12_reg[21]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__50_n_0));
  (* SOFT_HLUTNM = "soft_lutpair511" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__51
       (.I0(\TX_DATA_DEL12_reg[20]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__51_n_0));
  (* SOFT_HLUTNM = "soft_lutpair495" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__52
       (.I0(\TX_DATA_DEL12_reg[19]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__52_n_0));
  (* SOFT_HLUTNM = "soft_lutpair494" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__53
       (.I0(\TX_DATA_DEL12_reg[18]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__53_n_0));
  (* SOFT_HLUTNM = "soft_lutpair505" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__54
       (.I0(\TX_DATA_DEL12_reg[17]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__54_n_0));
  (* SOFT_HLUTNM = "soft_lutpair509" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__55
       (.I0(\TX_DATA_DEL12_reg[16]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__55_n_0));
  (* SOFT_HLUTNM = "soft_lutpair492" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__56
       (.I0(\TX_DATA_DEL12_reg[15]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__56_n_0));
  (* SOFT_HLUTNM = "soft_lutpair498" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__57
       (.I0(\TX_DATA_DEL12_reg[14]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__57_n_0));
  (* SOFT_HLUTNM = "soft_lutpair493" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__58
       (.I0(\TX_DATA_DEL12_reg[13]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__58_n_0));
  (* SOFT_HLUTNM = "soft_lutpair496" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__59
       (.I0(\TX_DATA_DEL12_reg[12]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__59_n_0));
  (* SOFT_HLUTNM = "soft_lutpair499" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__6
       (.I0(\TX_DATA_VALID_DEL12_reg[1]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair497" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__60
       (.I0(\TX_DATA_DEL12_reg[11]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__60_n_0));
  (* SOFT_HLUTNM = "soft_lutpair500" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__61
       (.I0(\TX_DATA_DEL12_reg[10]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__61_n_0));
  (* SOFT_HLUTNM = "soft_lutpair501" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__62
       (.I0(\TX_DATA_DEL12_reg[9]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__62_n_0));
  (* SOFT_HLUTNM = "soft_lutpair507" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__63
       (.I0(\TX_DATA_DEL12_reg[8]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__63_n_0));
  (* SOFT_HLUTNM = "soft_lutpair508" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__64
       (.I0(\TX_DATA_DEL12_reg[7]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__64_n_0));
  (* SOFT_HLUTNM = "soft_lutpair510" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__65
       (.I0(\TX_DATA_DEL12_reg[6]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__65_n_0));
  (* SOFT_HLUTNM = "soft_lutpair517" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__66
       (.I0(\TX_DATA_DEL12_reg[5]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__66_n_0));
  (* SOFT_HLUTNM = "soft_lutpair519" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__67
       (.I0(\TX_DATA_DEL12_reg[4]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__67_n_0));
  (* SOFT_HLUTNM = "soft_lutpair520" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__68
       (.I0(\TX_DATA_DEL12_reg[3]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__68_n_0));
  (* SOFT_HLUTNM = "soft_lutpair521" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__69
       (.I0(\TX_DATA_DEL12_reg[2]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__69_n_0));
  (* SOFT_HLUTNM = "soft_lutpair500" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__7
       (.I0(\TX_DATA_VALID_DEL12_reg[0]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair522" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__70
       (.I0(\TX_DATA_DEL12_reg[1]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__70_n_0));
  (* SOFT_HLUTNM = "soft_lutpair523" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__71
       (.I0(\TX_DATA_DEL12_reg[0]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__71_n_0));
  (* SOFT_HLUTNM = "soft_lutpair501" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__8
       (.I0(\TX_DATA_DEL12_reg[63]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__8_n_0));
  (* SOFT_HLUTNM = "soft_lutpair502" *) 
  LUT2 #(
    .INIT(4'h8)) 
    activity_blocks_gate__9
       (.I0(\TX_DATA_DEL12_reg[62]_activity_blocks_c_8_n_0 ),
        .I1(load_final_CRC_reg_0),
        .O(activity_blocks_gate__9_n_0));
  FDCE #(
    .INIT(1'b0)) 
    append_end_frame_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(txstatplus_int0_out[1]),
        .Q(append_end_frame));
  (* srl_bus_name = "\activity_blocks[0].dutH/append_reg_reg " *) 
  (* srl_name = "\activity_blocks[0].dutH/append_reg_reg[8]_srl9_activity_blocks_c_7 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \append_reg_reg[8]_srl9_activity_blocks_c_7 
       (.A0(1'b0),
        .A1(1'b0),
        .A2(1'b0),
        .A3(1'b1),
        .CE(1'b1),
        .CLK(clk_i),
        .D(load_CRC8),
        .Q(\append_reg_reg[8]_srl9_activity_blocks_c_7_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \append_reg_reg[9]_activity_blocks_c_8 
       (.C(clk_i),
        .CE(1'b1),
        .D(\append_reg_reg[8]_srl9_activity_blocks_c_7_n_0 ),
        .Q(\append_reg_reg[9]_activity_blocks_c_8_n_0 ),
        .R(1'b0));
  (* SOFT_HLUTNM = "soft_lutpair515" *) 
  LUT2 #(
    .INIT(4'h2)) 
    append_start_pause_i_1
       (.I0(transmit_pause_frame_reg_n_0),
        .I1(transmit_pause_frame_del),
        .O(append_start_pause0));
  FDCE #(
    .INIT(1'b0)) 
    append_start_pause_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(append_start_pause0),
        .Q(append_start_pause));
  FDCE #(
    .INIT(1'b0)) 
    apply_pause_delay_reg
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(apply_pause_delay),
        .Q(apply_pause_delay_reg_n_0));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[10]),
        .Q(byte_count_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[11]),
        .Q(byte_count_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[12]),
        .Q(byte_count_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[13]),
        .Q(byte_count_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[14]),
        .Q(byte_count_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[15]),
        .Q(byte_count_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[2]),
        .Q(byte_count_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[3]),
        .Q(byte_count_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[4]),
        .Q(byte_count_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[5]),
        .Q(byte_count_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[6]),
        .Q(byte_count_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[7]),
        .Q(byte_count_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[8]),
        .Q(byte_count_reg[8]));
  FDCE #(
    .INIT(1'b0)) 
    \byte_count_reg_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(BYTE_COUNTER[9]),
        .Q(byte_count_reg[9]));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[0]),
        .Q(\byte_count_stat_reg_n_0_[0] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[10]),
        .Q(\byte_count_stat_reg_n_0_[10] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[11]),
        .Q(\byte_count_stat_reg_n_0_[11] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[12]),
        .Q(\byte_count_stat_reg_n_0_[12] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[13]),
        .Q(\byte_count_stat_reg_n_0_[13] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[1]),
        .Q(\byte_count_stat_reg_n_0_[1] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[2]),
        .Q(\byte_count_stat_reg_n_0_[2] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[3]),
        .Q(\byte_count_stat_reg_n_0_[3] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[4]),
        .Q(\byte_count_stat_reg_n_0_[4] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[5]),
        .Q(\byte_count_stat_reg_n_0_[5] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[6]),
        .Q(\byte_count_stat_reg_n_0_[6] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[7]),
        .Q(\byte_count_stat_reg_n_0_[7] ),
        .R(transmit_pause_frame_reg_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \byte_count_stat_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[8]),
        .Q(\byte_count_stat_reg_n_0_[8] ),
        .R(transmit_pause_frame_reg_n_0));
  FDSE #(
    .INIT(1'b1)) 
    \byte_count_stat_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(final_byte_count_reg[9]),
        .Q(\byte_count_stat_reg_n_0_[9] ),
        .S(transmit_pause_frame_reg_n_0));
  FDPE #(
    .INIT(1'b1)) 
    fcs_enabled_int_reg
       (.C(clk_i),
        .CE(TX_CFG_REG_VALID),
        .D(TX_CFG_REG_VALUE[2]),
        .PRE(rst_i),
        .Q(fcs_enabled_int));
  LUT2 #(
    .INIT(4'h1)) 
    \final_byte_count[0]_i_1 
       (.I0(load_CRC8),
        .I1(final_byte_count_reg[0]),
        .O(p_0_in__2[0]));
  (* SOFT_HLUTNM = "soft_lutpair426" *) 
  LUT5 #(
    .INIT(32'hDFFFFFFF)) 
    \final_byte_count[10]_i_2 
       (.I0(final_byte_count_reg[8]),
        .I1(\final_byte_count[7]_i_2_n_0 ),
        .I2(final_byte_count_reg[6]),
        .I3(final_byte_count_reg[7]),
        .I4(final_byte_count_reg[9]),
        .O(\final_byte_count[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \final_byte_count[12]_i_2 
       (.I0(final_byte_count_reg[9]),
        .I1(final_byte_count_reg[7]),
        .I2(final_byte_count_reg[6]),
        .I3(\final_byte_count[7]_i_2_n_0 ),
        .I4(final_byte_count_reg[8]),
        .I5(final_byte_count_reg[10]),
        .O(\final_byte_count[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \final_byte_count[13]_i_2 
       (.I0(final_byte_count_reg[11]),
        .I1(final_byte_count_reg[10]),
        .I2(final_byte_count_reg[8]),
        .I3(\final_byte_count[7]_i_2_n_0 ),
        .I4(\final_byte_count[13]_i_3_n_0 ),
        .I5(final_byte_count_reg[9]),
        .O(\final_byte_count[13]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair490" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \final_byte_count[13]_i_3 
       (.I0(final_byte_count_reg[7]),
        .I1(final_byte_count_reg[6]),
        .O(\final_byte_count[13]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \final_byte_count[15]_i_3 
       (.I0(final_byte_count_reg[13]),
        .I1(final_byte_count_reg[11]),
        .I2(\final_byte_count[12]_i_2_n_0 ),
        .I3(final_byte_count_reg[12]),
        .O(\final_byte_count[15]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair491" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \final_byte_count[1]_i_1 
       (.I0(final_byte_count_reg[1]),
        .I1(final_byte_count_reg[0]),
        .I2(load_CRC8),
        .O(p_0_in__2[1]));
  (* SOFT_HLUTNM = "soft_lutpair491" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \final_byte_count[3]_i_2 
       (.I0(final_byte_count_reg[1]),
        .I1(final_byte_count_reg[0]),
        .I2(final_byte_count_reg[2]),
        .O(\final_byte_count[3]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair428" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \final_byte_count[4]_i_2 
       (.I0(final_byte_count_reg[2]),
        .I1(final_byte_count_reg[0]),
        .I2(final_byte_count_reg[1]),
        .I3(final_byte_count_reg[3]),
        .O(\final_byte_count[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair428" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \final_byte_count[5]_i_3 
       (.I0(final_byte_count_reg[3]),
        .I1(final_byte_count_reg[1]),
        .I2(final_byte_count_reg[0]),
        .I3(final_byte_count_reg[2]),
        .I4(final_byte_count_reg[4]),
        .O(\final_byte_count[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \final_byte_count[7]_i_2 
       (.I0(final_byte_count_reg[4]),
        .I1(final_byte_count_reg[2]),
        .I2(final_byte_count_reg[0]),
        .I3(final_byte_count_reg[1]),
        .I4(final_byte_count_reg[3]),
        .I5(final_byte_count_reg[5]),
        .O(\final_byte_count[7]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair490" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \final_byte_count[8]_i_2 
       (.I0(\final_byte_count[7]_i_2_n_0 ),
        .I1(final_byte_count_reg[6]),
        .I2(final_byte_count_reg[7]),
        .O(\final_byte_count[8]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair426" *) 
  LUT4 #(
    .INIT(16'hF7FF)) 
    \final_byte_count[9]_i_2 
       (.I0(final_byte_count_reg[7]),
        .I1(final_byte_count_reg[6]),
        .I2(\final_byte_count[7]_i_2_n_0 ),
        .I3(final_byte_count_reg[8]),
        .O(\final_byte_count[9]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[0] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[0]),
        .Q(final_byte_count_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[10] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[10]),
        .Q(final_byte_count_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[11] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[11]),
        .Q(final_byte_count_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[12] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[12]),
        .Q(final_byte_count_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[13] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[13]),
        .Q(final_byte_count_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[14] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[14]),
        .Q(final_byte_count_reg__0[14]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[15] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[15]),
        .Q(final_byte_count_reg__0[15]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[1] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[1]),
        .Q(final_byte_count_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[2] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[2]),
        .Q(final_byte_count_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[3] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[3]),
        .Q(final_byte_count_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[4] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[4]),
        .Q(final_byte_count_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[5] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[5]),
        .Q(final_byte_count_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[6] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[6]),
        .Q(final_byte_count_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[7] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[7]),
        .Q(final_byte_count_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[8] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[8]),
        .Q(final_byte_count_reg[8]));
  FDCE #(
    .INIT(1'b0)) 
    \final_byte_count_reg[9] 
       (.C(clk_i),
        .CE(U_CRC8_n_24),
        .CLR(rst_i),
        .D(p_0_in__2[9]),
        .Q(final_byte_count_reg[9]));
  FDCE #(
    .INIT(1'b0)) 
    frame_start_del_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(FRAME_START),
        .Q(frame_start_del));
  LUT5 #(
    .INIT(32'h00070004)) 
    insert_error_i_1
       (.I0(insert_error_i_2_n_0),
        .I1(load_CRC8),
        .I2(append_end_frame),
        .I3(reset_err_pause),
        .I4(txstatplus_int),
        .O(insert_error_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    insert_error_i_10
       (.I0(length_register[7]),
        .I1(final_byte_count_reg[7]),
        .I2(final_byte_count_reg[12]),
        .I3(final_byte_count_reg[13]),
        .I4(final_byte_count_reg[8]),
        .I5(final_byte_count_reg[9]),
        .O(insert_error_i_10_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    insert_error_i_11
       (.I0(final_byte_count_reg__0[14]),
        .I1(length_register[14]),
        .I2(final_byte_count_reg[11]),
        .I3(final_byte_count_reg[10]),
        .O(insert_error_i_11_n_0));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    insert_error_i_12
       (.I0(final_byte_count_reg[13]),
        .I1(length_register[13]),
        .I2(final_byte_count_reg[12]),
        .I3(length_register[12]),
        .I4(final_byte_count_reg__0[14]),
        .I5(length_register[14]),
        .O(insert_error_i_12_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    insert_error_i_13
       (.I0(final_byte_count_reg[6]),
        .I1(length_register[6]),
        .I2(final_byte_count_reg[8]),
        .I3(length_register[8]),
        .I4(final_byte_count_reg[7]),
        .I5(length_register[7]),
        .O(insert_error_i_13_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    insert_error_i_14
       (.I0(length_register[9]),
        .I1(final_byte_count_reg[9]),
        .I2(final_byte_count_reg[11]),
        .I3(length_register[11]),
        .I4(final_byte_count_reg[10]),
        .I5(length_register[10]),
        .O(insert_error_i_14_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    insert_error_i_15
       (.I0(length_register[0]),
        .I1(final_byte_count_reg[0]),
        .I2(final_byte_count_reg[2]),
        .I3(length_register[2]),
        .I4(final_byte_count_reg[1]),
        .I5(length_register[1]),
        .O(insert_error_i_15_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    insert_error_i_16
       (.I0(length_register[3]),
        .I1(final_byte_count_reg[3]),
        .I2(final_byte_count_reg[4]),
        .I3(length_register[4]),
        .I4(final_byte_count_reg[5]),
        .I5(length_register[5]),
        .O(insert_error_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair445" *) 
  LUT2 #(
    .INIT(4'h6)) 
    insert_error_i_17
       (.I0(final_byte_count_reg__0[15]),
        .I1(length_register[15]),
        .O(insert_error_i_17_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    insert_error_i_18
       (.I0(final_byte_count_reg[10]),
        .I1(final_byte_count_reg[11]),
        .O(insert_error_i_18_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    insert_error_i_19
       (.I0(final_byte_count_reg[8]),
        .I1(final_byte_count_reg[9]),
        .O(insert_error_i_19_n_0));
  LUT6 #(
    .INIT(64'h00000000FF040004)) 
    insert_error_i_2
       (.I0(insert_error_i_3_n_0),
        .I1(insert_error_i_4_n_0),
        .I2(insert_error_i_5_n_0),
        .I3(insert_error_i_6_n_0),
        .I4(insert_error1__0),
        .I5(tx_undderrun_int),
        .O(insert_error_i_2_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    insert_error_i_20
       (.I0(final_byte_count_reg[6]),
        .I1(final_byte_count_reg[7]),
        .O(insert_error_i_20_n_0));
  LUT3 #(
    .INIT(8'h4F)) 
    insert_error_i_21
       (.I0(final_byte_count_reg[4]),
        .I1(MAX_FRAME_SIZE[4]),
        .I2(final_byte_count_reg[5]),
        .O(insert_error_i_21_n_0));
  LUT4 #(
    .INIT(16'h44D4)) 
    insert_error_i_22
       (.I0(final_byte_count_reg[3]),
        .I1(MAX_FRAME_SIZE[3]),
        .I2(MAX_FRAME_SIZE[2]),
        .I3(final_byte_count_reg[2]),
        .O(insert_error_i_22_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    insert_error_i_23
       (.I0(final_byte_count_reg[1]),
        .O(insert_error_i_23_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    insert_error_i_24
       (.I0(final_byte_count_reg__0[15]),
        .I1(final_byte_count_reg__0[14]),
        .O(insert_error_i_24_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    insert_error_i_25
       (.I0(final_byte_count_reg[12]),
        .I1(final_byte_count_reg[13]),
        .O(insert_error_i_25_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    insert_error_i_26
       (.I0(final_byte_count_reg[10]),
        .I1(final_byte_count_reg[11]),
        .O(insert_error_i_26_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    insert_error_i_27
       (.I0(final_byte_count_reg[8]),
        .I1(final_byte_count_reg[9]),
        .O(insert_error_i_27_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    insert_error_i_28
       (.I0(final_byte_count_reg[7]),
        .I1(final_byte_count_reg[6]),
        .O(insert_error_i_28_n_0));
  LUT3 #(
    .INIT(8'h82)) 
    insert_error_i_29
       (.I0(final_byte_count_reg[5]),
        .I1(MAX_FRAME_SIZE[4]),
        .I2(final_byte_count_reg[4]),
        .O(insert_error_i_29_n_0));
  LUT5 #(
    .INIT(32'hFFFF8000)) 
    insert_error_i_3
       (.I0(length_register[4]),
        .I1(length_register[3]),
        .I2(length_register[5]),
        .I3(length_register[2]),
        .I4(insert_error_i_8_n_0),
        .O(insert_error_i_3_n_0));
  LUT4 #(
    .INIT(16'h9009)) 
    insert_error_i_30
       (.I0(MAX_FRAME_SIZE[3]),
        .I1(final_byte_count_reg[3]),
        .I2(MAX_FRAME_SIZE[2]),
        .I3(final_byte_count_reg[2]),
        .O(insert_error_i_30_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    insert_error_i_31
       (.I0(final_byte_count_reg[1]),
        .I1(final_byte_count_reg[0]),
        .O(insert_error_i_31_n_0));
  LUT5 #(
    .INIT(32'h00000010)) 
    insert_error_i_4
       (.I0(final_byte_count_reg[5]),
        .I1(length_register[9]),
        .I2(final_byte_count_reg[6]),
        .I3(length_register[6]),
        .I4(insert_error_i_9_n_0),
        .O(insert_error_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    insert_error_i_5
       (.I0(insert_error_i_10_n_0),
        .I1(insert_error_i_11_n_0),
        .I2(final_byte_count_reg[1]),
        .I3(final_byte_count_reg[0]),
        .I4(length_register[13]),
        .I5(length_register[15]),
        .O(insert_error_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    insert_error_i_6
       (.I0(insert_error_i_12_n_0),
        .I1(insert_error_i_13_n_0),
        .I2(insert_error_i_14_n_0),
        .I3(insert_error_i_15_n_0),
        .I4(insert_error_i_16_n_0),
        .I5(insert_error_i_17_n_0),
        .O(insert_error_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair445" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    insert_error_i_8
       (.I0(length_register[10]),
        .I1(final_byte_count_reg__0[15]),
        .I2(length_register[8]),
        .I3(final_byte_count_reg[4]),
        .O(insert_error_i_8_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    insert_error_i_9
       (.I0(length_register[12]),
        .I1(final_byte_count_reg[3]),
        .I2(length_register[11]),
        .I3(final_byte_count_reg[2]),
        .O(insert_error_i_9_n_0));
  FDCE #(
    .INIT(1'b0)) 
    insert_error_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(insert_error_i_1_n_0),
        .Q(txstatplus_int));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    insert_error_reg_i_7
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({insert_error1__0,insert_error_reg_i_7_n_1,insert_error_reg_i_7_n_2,insert_error_reg_i_7_n_3,insert_error_reg_i_7_n_4,insert_error_reg_i_7_n_5,insert_error_reg_i_7_n_6,insert_error_reg_i_7_n_7}),
        .DI({1'b0,1'b0,insert_error_i_18_n_0,insert_error_i_19_n_0,insert_error_i_20_n_0,insert_error_i_21_n_0,insert_error_i_22_n_0,insert_error_i_23_n_0}),
        .O(NLW_insert_error_reg_i_7_O_UNCONNECTED[7:0]),
        .S({insert_error_i_24_n_0,insert_error_i_25_n_0,insert_error_i_26_n_0,insert_error_i_27_n_0,insert_error_i_28_n_0,insert_error_i_29_n_0,insert_error_i_30_n_0,insert_error_i_31_n_0}));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[0] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_43),
        .Q(length_register[0]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[10] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_33),
        .Q(length_register[10]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[11] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_32),
        .Q(length_register[11]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[12] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_31),
        .Q(length_register[12]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[13] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_30),
        .Q(length_register[13]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[14] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_29),
        .Q(length_register[14]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[15] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_28),
        .Q(length_register[15]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[1] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_42),
        .Q(length_register[1]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[2] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_41),
        .Q(length_register[2]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[3] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_40),
        .Q(length_register[3]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[4] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_39),
        .Q(length_register[4]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[5] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_38),
        .Q(length_register[5]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[6] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_37),
        .Q(length_register[6]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[7] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_36),
        .Q(length_register[7]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[8] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_35),
        .Q(length_register[8]));
  FDCE #(
    .INIT(1'b0)) 
    \length_register_reg[9] 
       (.C(clk_i),
        .CE(length_register0),
        .CLR(rst_i),
        .D(U_byte_count_module_n_34),
        .Q(length_register[9]));
  LUT4 #(
    .INIT(16'h4F44)) 
    load_CRC8_i_1
       (.I0(transmit_pause_frame_del2),
        .I1(transmit_pause_frame_del3),
        .I2(FRAME_START),
        .I3(frame_start_del),
        .O(load_CRC80));
  FDCE #(
    .INIT(1'b0)) 
    load_CRC8_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(load_CRC80),
        .Q(load_CRC8));
  FDCE #(
    .INIT(1'b0)) 
    load_final_CRC_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(activity_blocks_gate_n_0),
        .Q(txstatplus_int0_out[1]));
  (* SOFT_HLUTNM = "soft_lutpair506" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \pause_frame_counter[0]_i_1 
       (.I0(pause_frame_counter_reg[0]),
        .O(\pause_frame_counter[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair506" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \pause_frame_counter[1]_i_1 
       (.I0(pause_frame_counter_reg[0]),
        .I1(pause_frame_counter_reg[1]),
        .O(p_0_in__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair440" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \pause_frame_counter[2]_i_1 
       (.I0(pause_frame_counter_reg[2]),
        .I1(pause_frame_counter_reg[1]),
        .I2(pause_frame_counter_reg[0]),
        .O(p_0_in__0[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \pause_frame_counter[3]_i_1 
       (.I0(transmit_pause_frame_reg_n_0),
        .I1(FRAME_START),
        .O(pause_frame_counter0));
  (* SOFT_HLUTNM = "soft_lutpair440" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \pause_frame_counter[3]_i_2 
       (.I0(pause_frame_counter_reg[3]),
        .I1(pause_frame_counter_reg[0]),
        .I2(pause_frame_counter_reg[1]),
        .I3(pause_frame_counter_reg[2]),
        .O(p_0_in__0[3]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_counter_reg[0] 
       (.C(clk_i),
        .CE(pause_frame_counter0),
        .CLR(rst_i),
        .D(\pause_frame_counter[0]_i_1_n_0 ),
        .Q(pause_frame_counter_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_counter_reg[1] 
       (.C(clk_i),
        .CE(pause_frame_counter0),
        .CLR(rst_i),
        .D(p_0_in__0[1]),
        .Q(pause_frame_counter_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_counter_reg[2] 
       (.C(clk_i),
        .CE(pause_frame_counter0),
        .CLR(rst_i),
        .D(p_0_in__0[2]),
        .Q(pause_frame_counter_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_counter_reg[3] 
       (.C(clk_i),
        .CE(pause_frame_counter0),
        .CLR(rst_i),
        .D(p_0_in__0[3]),
        .Q(pause_frame_counter_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    read_ifg_int_reg
       (.C(clk_i),
        .CE(TX_CFG_REG_VALID),
        .CLR(rst_i),
        .D(TX_CFG_REG_VALUE[0]),
        .Q(read_ifg_int));
  (* SOFT_HLUTNM = "soft_lutpair515" *) 
  LUT2 #(
    .INIT(4'h2)) 
    reset_err_pause_i_1
       (.I0(transmit_pause_frame_del),
        .I1(transmit_pause_frame_reg_n_0),
        .O(reset_err_pause0));
  FDCE #(
    .INIT(1'b0)) 
    reset_err_pause_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(reset_err_pause0),
        .Q(reset_err_pause));
  FDCE #(
    .INIT(1'b0)) 
    reset_tx_int_reg
       (.C(clk_i),
        .CE(TX_CFG_REG_VALID),
        .CLR(rst_i),
        .D(TX_CFG_REG_VALUE[3]),
        .Q(reset_tx_int));
  LUT1 #(
    .INIT(2'h1)) 
    \rp[1]_i_3 
       (.I0(rst_i),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair487" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    set_pause_stats_i_1
       (.I0(PAUSEVAL_DEL2),
        .I1(append_end_frame),
        .I2(set_pause_stats),
        .O(set_pause_stats_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    set_pause_stats_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(set_pause_stats_i_1_n_0),
        .Q(set_pause_stats));
  LUT6 #(
    .INIT(64'h00000E0000000200)) 
    \shift_pause_data[0]_i_1 
       (.I0(TXD_PAUSE_DEL1),
        .I1(pause_frame_counter_reg[0]),
        .I2(pause_frame_counter_reg[1]),
        .I3(\shift_pause_valid[0]_i_1_n_0 ),
        .I4(pause_frame_counter_reg[2]),
        .I5(TXD_PAUSE_DEL2[0]),
        .O(\shift_pause_data[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair535" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[10]_i_1 
       (.I0(TXD_PAUSE_DEL2[10]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair534" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[11]_i_1 
       (.I0(TXD_PAUSE_DEL2[11]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair533" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[12]_i_1 
       (.I0(TXD_PAUSE_DEL2[12]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair532" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[13]_i_1 
       (.I0(TXD_PAUSE_DEL2[13]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair531" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[14]_i_1 
       (.I0(TXD_PAUSE_DEL2[14]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair530" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[15]_i_1 
       (.I0(TXD_PAUSE_DEL2[15]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair529" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[1]_i_1 
       (.I0(TXD_PAUSE_DEL2[1]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair530" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[2]_i_1 
       (.I0(TXD_PAUSE_DEL2[2]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair531" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[3]_i_1 
       (.I0(TXD_PAUSE_DEL2[3]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair532" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[4]_i_1 
       (.I0(TXD_PAUSE_DEL2[4]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair529" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[56]_i_1 
       (.I0(TXD_PAUSE_DEL1),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[56]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    \shift_pause_data[56]_i_2 
       (.I0(pause_frame_counter_reg[0]),
        .I1(pause_frame_counter_reg[1]),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_reg_n_0),
        .I4(pause_frame_counter_reg[3]),
        .I5(pause_frame_counter_reg[2]),
        .O(\shift_pause_data[56]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair533" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[5]_i_1 
       (.I0(TXD_PAUSE_DEL2[5]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \shift_pause_data[60]_i_1 
       (.I0(pause_frame_counter_reg[0]),
        .I1(pause_frame_counter_reg[1]),
        .I2(TXD_PAUSE_DEL1),
        .I3(pause_frame_counter0),
        .I4(pause_frame_counter_reg[3]),
        .I5(pause_frame_counter_reg[2]),
        .O(\shift_pause_data[60]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair534" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[6]_i_1 
       (.I0(TXD_PAUSE_DEL2[6]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair535" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[7]_i_1 
       (.I0(TXD_PAUSE_DEL2[7]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000E0000000200)) 
    \shift_pause_data[8]_i_1 
       (.I0(TXD_PAUSE_DEL1),
        .I1(pause_frame_counter_reg[0]),
        .I2(pause_frame_counter_reg[1]),
        .I3(\shift_pause_valid[0]_i_1_n_0 ),
        .I4(pause_frame_counter_reg[2]),
        .I5(TXD_PAUSE_DEL2[8]),
        .O(\shift_pause_data[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \shift_pause_data[9]_i_1 
       (.I0(TXD_PAUSE_DEL2[9]),
        .I1(\shift_pause_data[56]_i_2_n_0 ),
        .O(\shift_pause_data[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[0]_i_1_n_0 ),
        .Q(shift_pause_data[0]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[10]_i_1_n_0 ),
        .Q(shift_pause_data[10]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[11]_i_1_n_0 ),
        .Q(shift_pause_data[11]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[12]_i_1_n_0 ),
        .Q(shift_pause_data[12]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[13]_i_1_n_0 ),
        .Q(shift_pause_data[13]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[14]_i_1_n_0 ),
        .Q(shift_pause_data[14]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[15]_i_1_n_0 ),
        .Q(shift_pause_data[15]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[1]_i_1_n_0 ),
        .Q(shift_pause_data[1]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[2]_i_1_n_0 ),
        .Q(shift_pause_data[2]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[3]_i_1_n_0 ),
        .Q(shift_pause_data[3]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[4]_i_1_n_0 ),
        .Q(shift_pause_data[4]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[56]_i_1_n_0 ),
        .Q(shift_pause_data[56]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[5]_i_1_n_0 ),
        .Q(shift_pause_data[5]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[60]_i_1_n_0 ),
        .Q(shift_pause_data[60]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[6]_i_1_n_0 ),
        .Q(shift_pause_data[6]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[7]_i_1_n_0 ),
        .Q(shift_pause_data[7]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[8]_i_1_n_0 ),
        .Q(shift_pause_data[8]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_data_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_data[9]_i_1_n_0 ),
        .Q(shift_pause_data[9]));
  (* SOFT_HLUTNM = "soft_lutpair469" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \shift_pause_valid[0]_i_1 
       (.I0(FRAME_START),
        .I1(transmit_pause_frame_reg_n_0),
        .I2(pause_frame_counter_reg[3]),
        .O(\shift_pause_valid[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0004040404040404)) 
    \shift_pause_valid[4]_i_1 
       (.I0(pause_frame_counter_reg[3]),
        .I1(transmit_pause_frame_reg_n_0),
        .I2(FRAME_START),
        .I3(pause_frame_counter_reg[0]),
        .I4(pause_frame_counter_reg[1]),
        .I5(pause_frame_counter_reg[2]),
        .O(\shift_pause_valid[4]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_valid_del_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(shift_pause_valid[0]),
        .Q(shift_pause_valid_del[0]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_valid_del_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(shift_pause_valid[4]),
        .Q(shift_pause_valid_del[4]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_valid_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_valid[0]_i_1_n_0 ),
        .Q(shift_pause_valid[0]));
  FDCE #(
    .INIT(1'b0)) 
    \shift_pause_valid_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\shift_pause_valid[4]_i_1_n_0 ),
        .Q(shift_pause_valid[4]));
  FDCE #(
    .INIT(1'b0)) 
    start_CRC8_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid_reg_n_0_[0] ),
        .Q(start_CRC8));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[0] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_39),
        .Q(store_pause_frame[0]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[10] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_29),
        .Q(store_pause_frame[10]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[11] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_28),
        .Q(store_pause_frame[11]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[12] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_27),
        .Q(store_pause_frame[12]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[13] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_26),
        .Q(store_pause_frame[13]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[14] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_25),
        .Q(store_pause_frame[14]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[15] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_24),
        .Q(store_pause_frame[15]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[1] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_38),
        .Q(store_pause_frame[1]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[2] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_37),
        .Q(store_pause_frame[2]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[3] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_36),
        .Q(store_pause_frame[3]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[4] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_35),
        .Q(store_pause_frame[4]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[5] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_34),
        .Q(store_pause_frame[5]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[6] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_33),
        .Q(store_pause_frame[6]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[7] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_32),
        .Q(store_pause_frame[7]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[8] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_31),
        .Q(store_pause_frame[8]));
  FDCE #(
    .INIT(1'b0)) 
    \store_pause_frame_reg[9] 
       (.C(clk_i),
        .CE(U_ACK_CNT_n_13),
        .CLR(rst_i),
        .D(U_ACK_CNT_n_30),
        .Q(store_pause_frame[9]));
  (* SOFT_HLUTNM = "soft_lutpair454" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[0]_i_1 
       (.I0(TX_DATA_DEL2[0]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[8] ),
        .O(\store_tx_data[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair464" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[10]_i_1 
       (.I0(TX_DATA_DEL2[10]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[18] ),
        .O(\store_tx_data[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair465" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[11]_i_1 
       (.I0(TX_DATA_DEL2[11]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[19] ),
        .O(\store_tx_data[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair466" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[12]_i_1 
       (.I0(TX_DATA_DEL2[12]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[20] ),
        .O(\store_tx_data[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair467" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[13]_i_1 
       (.I0(TX_DATA_DEL2[13]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[21] ),
        .O(\store_tx_data[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair468" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[14]_i_1 
       (.I0(TX_DATA_DEL2[14]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[22] ),
        .O(\store_tx_data[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair471" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[15]_i_1 
       (.I0(TX_DATA_DEL2[15]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[23] ),
        .O(\store_tx_data[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair472" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[16]_i_1 
       (.I0(TX_DATA_DEL2[16]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[24] ),
        .O(\store_tx_data[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair473" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[17]_i_1 
       (.I0(TX_DATA_DEL2[17]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[25] ),
        .O(\store_tx_data[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair474" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[18]_i_1 
       (.I0(TX_DATA_DEL2[18]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[26] ),
        .O(\store_tx_data[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair475" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[19]_i_1 
       (.I0(TX_DATA_DEL2[19]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[27] ),
        .O(\store_tx_data[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair455" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[1]_i_1 
       (.I0(TX_DATA_DEL2[1]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[9] ),
        .O(\store_tx_data[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair476" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[20]_i_1 
       (.I0(TX_DATA_DEL2[20]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[28] ),
        .O(\store_tx_data[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair477" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[21]_i_1 
       (.I0(TX_DATA_DEL2[21]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[29] ),
        .O(\store_tx_data[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair478" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[22]_i_1 
       (.I0(TX_DATA_DEL2[22]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[30] ),
        .O(\store_tx_data[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair479" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[23]_i_1 
       (.I0(TX_DATA_DEL2[23]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[31] ),
        .O(\store_tx_data[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair480" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[24]_i_1 
       (.I0(TX_DATA_DEL2[24]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[32] ),
        .O(\store_tx_data[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair481" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[25]_i_1 
       (.I0(TX_DATA_DEL2[25]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[33] ),
        .O(\store_tx_data[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair482" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[26]_i_1 
       (.I0(TX_DATA_DEL2[26]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[34] ),
        .O(\store_tx_data[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair483" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[27]_i_1 
       (.I0(TX_DATA_DEL2[27]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[35] ),
        .O(\store_tx_data[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair484" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[28]_i_1 
       (.I0(TX_DATA_DEL2[28]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[36] ),
        .O(\store_tx_data[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair485" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[29]_i_1 
       (.I0(TX_DATA_DEL2[29]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[37] ),
        .O(\store_tx_data[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair456" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[2]_i_1 
       (.I0(TX_DATA_DEL2[2]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[10] ),
        .O(\store_tx_data[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair486" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[30]_i_1 
       (.I0(TX_DATA_DEL2[30]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[38] ),
        .O(\store_tx_data[30]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[31]_i_1 
       (.I0(TX_DATA_DEL2[31]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[39] ),
        .O(\store_tx_data[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair486" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[32]_i_1 
       (.I0(TX_DATA_DEL2[32]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[40] ),
        .O(\store_tx_data[32]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair485" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[33]_i_1 
       (.I0(TX_DATA_DEL2[33]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[41] ),
        .O(\store_tx_data[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair484" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[34]_i_1 
       (.I0(TX_DATA_DEL2[34]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[42] ),
        .O(\store_tx_data[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair483" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[35]_i_1 
       (.I0(TX_DATA_DEL2[35]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[43] ),
        .O(\store_tx_data[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair482" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[36]_i_1 
       (.I0(TX_DATA_DEL2[36]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[44] ),
        .O(\store_tx_data[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair481" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[37]_i_1 
       (.I0(TX_DATA_DEL2[37]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[45] ),
        .O(\store_tx_data[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair480" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[38]_i_1 
       (.I0(TX_DATA_DEL2[38]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[46] ),
        .O(\store_tx_data[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair479" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[39]_i_1 
       (.I0(TX_DATA_DEL2[39]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[47] ),
        .O(\store_tx_data[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair457" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[3]_i_1 
       (.I0(TX_DATA_DEL2[3]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[11] ),
        .O(\store_tx_data[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair478" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[40]_i_1 
       (.I0(TX_DATA_DEL2[40]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[48] ),
        .O(\store_tx_data[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair477" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[41]_i_1 
       (.I0(TX_DATA_DEL2[41]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[49] ),
        .O(\store_tx_data[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair476" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[42]_i_1 
       (.I0(TX_DATA_DEL2[42]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[50] ),
        .O(\store_tx_data[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair475" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[43]_i_1 
       (.I0(TX_DATA_DEL2[43]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[51] ),
        .O(\store_tx_data[43]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair474" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[44]_i_1 
       (.I0(TX_DATA_DEL2[44]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[52] ),
        .O(\store_tx_data[44]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair473" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[45]_i_1 
       (.I0(TX_DATA_DEL2[45]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[53] ),
        .O(\store_tx_data[45]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair472" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[46]_i_1 
       (.I0(TX_DATA_DEL2[46]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[54] ),
        .O(\store_tx_data[46]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair471" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[47]_i_1 
       (.I0(TX_DATA_DEL2[47]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[55] ),
        .O(\store_tx_data[47]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair468" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[48]_i_1 
       (.I0(TX_DATA_DEL2[48]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[56] ),
        .O(\store_tx_data[48]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair467" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[49]_i_1 
       (.I0(TX_DATA_DEL2[49]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[57] ),
        .O(\store_tx_data[49]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair458" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[4]_i_1 
       (.I0(TX_DATA_DEL2[4]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[12] ),
        .O(\store_tx_data[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair466" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[50]_i_1 
       (.I0(TX_DATA_DEL2[50]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[58] ),
        .O(\store_tx_data[50]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair465" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[51]_i_1 
       (.I0(TX_DATA_DEL2[51]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[59] ),
        .O(\store_tx_data[51]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair464" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[52]_i_1 
       (.I0(TX_DATA_DEL2[52]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[60] ),
        .O(\store_tx_data[52]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair463" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[53]_i_1 
       (.I0(TX_DATA_DEL2[53]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[61] ),
        .O(\store_tx_data[53]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair462" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[54]_i_1 
       (.I0(TX_DATA_DEL2[54]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[62] ),
        .O(\store_tx_data[54]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair461" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[55]_i_1 
       (.I0(TX_DATA_DEL2[55]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[63] ),
        .O(\store_tx_data[55]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair459" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[5]_i_1 
       (.I0(TX_DATA_DEL2[5]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[13] ),
        .O(\store_tx_data[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair460" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[6]_i_1 
       (.I0(TX_DATA_DEL2[6]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[14] ),
        .O(\store_tx_data[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair461" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[7]_i_1 
       (.I0(TX_DATA_DEL2[7]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[15] ),
        .O(\store_tx_data[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair462" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[8]_i_1 
       (.I0(TX_DATA_DEL2[8]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[16] ),
        .O(\store_tx_data[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair463" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data[9]_i_1 
       (.I0(TX_DATA_DEL2[9]),
        .I1(load_CRC8),
        .I2(\store_tx_data_reg_n_0_[17] ),
        .O(\store_tx_data[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[0]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[10]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[11]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[12]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[13]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[14]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[15]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[16]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[17]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[18]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[19]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[1]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[20]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[21]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[22]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[23]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[24]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[25]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[26]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[27]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[28]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[29]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[2]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[30]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[31]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[32]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[32] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[33]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[33] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[34]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[34] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[35]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[35] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[36]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[36] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[37]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[37] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[38]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[38] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[39]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[39] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[3]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[40]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[40] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[41]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[41] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[42]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[42] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[43]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[43] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[44]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[44] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[45]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[45] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[46]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[46] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[47]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[47] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[48]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[48] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[49]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[49] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[4]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[50]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[50] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[51]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[51] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[52]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[52] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[53]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[53] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[54]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[54] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[55]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[55] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[56] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[56]),
        .Q(\store_tx_data_reg_n_0_[56] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[57] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[57]),
        .Q(\store_tx_data_reg_n_0_[57] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[58] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[58]),
        .Q(\store_tx_data_reg_n_0_[58] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[59] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[59]),
        .Q(\store_tx_data_reg_n_0_[59] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[5]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[60] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[60]),
        .Q(\store_tx_data_reg_n_0_[60] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[61] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[61]),
        .Q(\store_tx_data_reg_n_0_[61] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[62] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[62]),
        .Q(\store_tx_data_reg_n_0_[62] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[63] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_DEL2[63]),
        .Q(\store_tx_data_reg_n_0_[63] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[6]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[7]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[8]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data[9]_i_1_n_0 ),
        .Q(\store_tx_data_reg_n_0_[9] ));
  (* SOFT_HLUTNM = "soft_lutpair460" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[0]_i_1 
       (.I0(TX_DATA_VALID_DEL2[0]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[1] ),
        .O(\store_tx_data_valid[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair459" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[1]_i_1 
       (.I0(TX_DATA_VALID_DEL2[1]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[2] ),
        .O(\store_tx_data_valid[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair458" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[2]_i_1 
       (.I0(TX_DATA_VALID_DEL2[2]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[3] ),
        .O(\store_tx_data_valid[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair457" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[3]_i_1 
       (.I0(TX_DATA_VALID_DEL2[3]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[4] ),
        .O(\store_tx_data_valid[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair456" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[4]_i_1 
       (.I0(TX_DATA_VALID_DEL2[4]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[5] ),
        .O(\store_tx_data_valid[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair455" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[5]_i_1 
       (.I0(TX_DATA_VALID_DEL2[5]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[6] ),
        .O(\store_tx_data_valid[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair454" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \store_tx_data_valid[6]_i_1 
       (.I0(TX_DATA_VALID_DEL2[6]),
        .I1(load_CRC8),
        .I2(\store_tx_data_valid_reg_n_0_[7] ),
        .O(\store_tx_data_valid[6]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[0]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[1]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[2]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[3]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[4]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[5]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\store_tx_data_valid[6]_i_1_n_0 ),
        .Q(\store_tx_data_valid_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \store_tx_data_valid_reg[7] 
       (.C(clk_i),
        .CE(load_CRC8),
        .CLR(rst_i),
        .D(TX_DATA_VALID_DEL2[7]),
        .Q(\store_tx_data_valid_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    transmit_pause_frame_del2_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(transmit_pause_frame_del),
        .Q(transmit_pause_frame_del2));
  FDCE #(
    .INIT(1'b0)) 
    transmit_pause_frame_del3_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(transmit_pause_frame_del2),
        .Q(transmit_pause_frame_del3));
  FDCE #(
    .INIT(1'b0)) 
    transmit_pause_frame_del_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(transmit_pause_frame_reg_n_0),
        .Q(transmit_pause_frame_del));
  LUT6 #(
    .INIT(64'hFFFFFFEFAAAAAAAA)) 
    transmit_pause_frame_i_1
       (.I0(PAUSEVAL_DEL2),
        .I1(pause_frame_counter_reg[2]),
        .I2(pause_frame_counter_reg[3]),
        .I3(pause_frame_counter_reg[0]),
        .I4(pause_frame_counter_reg[1]),
        .I5(transmit_pause_frame_reg_n_0),
        .O(transmit_pause_frame_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    transmit_pause_frame_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(transmit_pause_frame_i_1_n_0),
        .Q(transmit_pause_frame_reg_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    transmit_pause_frame_valid_i_1
       (.I0(transmit_pause_frame_reg_n_0),
        .I1(transmit_pause_frame_del),
        .O(transmit_pause_frame_valid0));
  FDCE #(
    .INIT(1'b0)) 
    transmit_pause_frame_valid_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(transmit_pause_frame_valid0),
        .Q(transmit_pause_frame_valid));
  LUT1 #(
    .INIT(2'h1)) 
    \tx_data_int[7]_i_1 
       (.I0(load_CRC8),
        .O(\tx_data_int[7]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[0] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[0] ),
        .Q(tx_data_int[0]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[1] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[1] ),
        .Q(tx_data_int[1]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[2] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[2] ),
        .Q(tx_data_int[2]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[3] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[3] ),
        .Q(tx_data_int[3]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[4] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[4] ),
        .Q(tx_data_int[4]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[5] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[5] ),
        .Q(tx_data_int[5]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[6] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[6] ),
        .Q(tx_data_int[6]));
  FDCE #(
    .INIT(1'b0)) 
    \tx_data_int_reg[7] 
       (.C(clk_i),
        .CE(\tx_data_int[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\store_tx_data_reg_n_0_[7] ),
        .Q(tx_data_int[7]));
  LUT4 #(
    .INIT(16'h0054)) 
    tx_undderrun_int_i_1
       (.I0(rst_i),
        .I1(tx_undderrun_int_reg_0),
        .I2(tx_undderrun_int),
        .I3(append_end_frame),
        .O(tx_undderrun_int_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    tx_undderrun_int_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(tx_undderrun_int_i_1_n_0),
        .Q(tx_undderrun_int),
        .R(1'b0));
  (* SOFT_HLUTNM = "soft_lutpair438" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[10]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[5] ),
        .O(txstatplus_int0_out[10]));
  (* SOFT_HLUTNM = "soft_lutpair439" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[11]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[6] ),
        .O(txstatplus_int0_out[11]));
  (* SOFT_HLUTNM = "soft_lutpair439" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[12]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[7] ),
        .O(txstatplus_int0_out[12]));
  (* SOFT_HLUTNM = "soft_lutpair438" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[13]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[8] ),
        .O(txstatplus_int0_out[13]));
  (* SOFT_HLUTNM = "soft_lutpair437" *) 
  LUT4 #(
    .INIT(16'hAAA8)) 
    \txstatplus_int[14]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(final_byte_count_reg__0[15]),
        .I2(\byte_count_stat_reg_n_0_[9] ),
        .I3(vlan_enabled_int),
        .O(txstatplus_int0_out[14]));
  (* SOFT_HLUTNM = "soft_lutpair436" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[15]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[10] ),
        .O(txstatplus_int0_out[15]));
  (* SOFT_HLUTNM = "soft_lutpair435" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[16]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[11] ),
        .O(txstatplus_int0_out[16]));
  (* SOFT_HLUTNM = "soft_lutpair434" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[17]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[12] ),
        .O(txstatplus_int0_out[17]));
  LUT3 #(
    .INIT(8'hDF)) 
    \txstatplus_int[18]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(set_pause_stats),
        .I2(vlan_enabled_int),
        .O(\txstatplus_int[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair433" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[18]_i_2 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[13] ),
        .O(txstatplus_int0_out[18]));
  (* SOFT_HLUTNM = "soft_lutpair446" *) 
  LUT3 #(
    .INIT(8'hC8)) 
    \txstatplus_int[19]_i_1 
       (.I0(vlan_enabled_int),
        .I1(txstatplus_int0_out[1]),
        .I2(\txstatplus_int_reg_n_0_[19] ),
        .O(\txstatplus_int[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \txstatplus_int[24]_i_1 
       (.I0(set_pause_stats),
        .I1(txstatplus_int0_out[1]),
        .O(\txstatplus_int[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair447" *) 
  LUT3 #(
    .INIT(8'hC8)) 
    \txstatplus_int[3]_i_1 
       (.I0(txstatplus_int),
        .I1(txstatplus_int0_out[1]),
        .I2(\txstatplus_int_reg_n_0_[3] ),
        .O(\txstatplus_int[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair433" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[5]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[0] ),
        .O(txstatplus_int0_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair434" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[6]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[1] ),
        .O(txstatplus_int0_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair435" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[7]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[2] ),
        .O(txstatplus_int0_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair436" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[8]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[3] ),
        .O(txstatplus_int0_out[8]));
  (* SOFT_HLUTNM = "soft_lutpair437" *) 
  LUT4 #(
    .INIT(16'h2220)) 
    \txstatplus_int[9]_i_1 
       (.I0(txstatplus_int0_out[1]),
        .I1(vlan_enabled_int),
        .I2(final_byte_count_reg__0[15]),
        .I3(\byte_count_stat_reg_n_0_[4] ),
        .O(txstatplus_int0_out[9]));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[10] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[10]),
        .Q(\txstatplus_int_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[11] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[11]),
        .Q(\txstatplus_int_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[12] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[12]),
        .Q(\txstatplus_int_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[13] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[13]),
        .Q(\txstatplus_int_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[14] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[14]),
        .Q(\txstatplus_int_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[15] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[15]),
        .Q(\txstatplus_int_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[16] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[16]),
        .Q(\txstatplus_int_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[17] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[17]),
        .Q(\txstatplus_int_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[18] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[18]),
        .Q(\txstatplus_int_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\txstatplus_int[19]_i_1_n_0 ),
        .Q(\txstatplus_int_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[1] 
       (.C(clk_i),
        .CE(\txstatplus_int[24]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[1]),
        .Q(\txstatplus_int_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[24] 
       (.C(clk_i),
        .CE(\txstatplus_int[24]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[1]),
        .Q(\txstatplus_int_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[2] 
       (.C(clk_i),
        .CE(\txstatplus_int[24]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[1]),
        .Q(\txstatplus_int_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\txstatplus_int[3]_i_1_n_0 ),
        .Q(\txstatplus_int_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[4] 
       (.C(clk_i),
        .CE(\txstatplus_int[24]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[1]),
        .Q(\txstatplus_int_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[5] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[5]),
        .Q(\txstatplus_int_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[6] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[6]),
        .Q(\txstatplus_int_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[7] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[7]),
        .Q(\txstatplus_int_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[8] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[8]),
        .Q(\txstatplus_int_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \txstatplus_int_reg[9] 
       (.C(clk_i),
        .CE(\txstatplus_int[18]_i_1_n_0 ),
        .CLR(rst_i),
        .D(txstatplus_int0_out[9]),
        .Q(\txstatplus_int_reg_n_0_[9] ));
  FDCE #(
    .INIT(1'b0)) 
    vlan_enabled_int_reg
       (.C(clk_i),
        .CE(TX_CFG_REG_VALID),
        .CLR(rst_i),
        .D(TX_CFG_REG_VALUE[1]),
        .Q(vlan_enabled_int));
endmodule

(* ORIG_REF_NAME = "ack_counter" *) 
module switch_elements_ack_counter
   (tx_ack_reg_0,
    D,
    append_start_pause_reg,
    append_start_pause_reg_0,
    E,
    apply_pause_delay,
    AR,
    tx_ack_reg_1,
    tx_ack_reg_2,
    tx_ack_reg_3,
    tx_ack_reg_4,
    tx_ack_reg_5,
    tx_ack_reg_6,
    tx_ack_reg_7,
    SS,
    \FC_TX_PAUSEDATA_reg[15] ,
    clk_i,
    out,
    rst_i,
    reset_tx_int,
    Q,
    \TX_DATA_REG_reg[63] ,
    \TX_DATA_REG_reg[63]_0 ,
    FRAME_START,
    \TX_DATA_REG_reg[63]_1 ,
    apply_pause_delay_reg,
    \TX_DATA_REG_reg[40] ,
    append_start_pause,
    transmit_pause_frame_valid,
    I94,
    start_count_del_reg_0);
  output tx_ack_reg_0;
  output [9:0]D;
  output append_start_pause_reg;
  output append_start_pause_reg_0;
  output [0:0]E;
  output apply_pause_delay;
  output [0:0]AR;
  output tx_ack_reg_1;
  output tx_ack_reg_2;
  output tx_ack_reg_3;
  output tx_ack_reg_4;
  output tx_ack_reg_5;
  output tx_ack_reg_6;
  output tx_ack_reg_7;
  output [0:0]SS;
  output [15:0]\FC_TX_PAUSEDATA_reg[15] ;
  input clk_i;
  input out;
  input rst_i;
  input reset_tx_int;
  input [15:0]Q;
  input \TX_DATA_REG_reg[63] ;
  input [1:0]\TX_DATA_REG_reg[63]_0 ;
  input FRAME_START;
  input [9:0]\TX_DATA_REG_reg[63]_1 ;
  input apply_pause_delay_reg;
  input [11:0]\TX_DATA_REG_reg[40] ;
  input append_start_pause;
  input transmit_pause_frame_valid;
  input [15:0]I94;
  input start_count_del_reg_0;

  wire [0:0]AR;
  wire [9:0]D;
  wire [0:0]E;
  wire [15:0]\FC_TX_PAUSEDATA_reg[15] ;
  wire FRAME_START;
  wire [15:0]I94;
  wire [15:0]Q;
  wire [0:0]SS;
  wire [11:0]\TX_DATA_REG_reg[40] ;
  wire \TX_DATA_REG_reg[63] ;
  wire [1:0]\TX_DATA_REG_reg[63]_0 ;
  wire [9:0]\TX_DATA_REG_reg[63]_1 ;
  wire append_start_pause;
  wire append_start_pause_reg;
  wire append_start_pause_reg_0;
  wire apply_pause_delay;
  wire apply_pause_delay_reg;
  wire clk_i;
  wire \counter[10]_i_2_n_0 ;
  wire \counter[14]_i_2_n_0 ;
  wire \counter[15]_i_1__0_n_0 ;
  wire \counter[15]_i_3_n_0 ;
  wire \counter[5]_i_2_n_0 ;
  wire \counter[9]_i_2_n_0 ;
  wire [15:0]counter_reg;
  wire out;
  wire [15:0]p_0_in;
  wire reset0;
  wire reset_tx_int;
  wire rst_i;
  wire start_count;
  wire start_count_del;
  wire start_count_del_reg_0;
  wire start_count_reg_i_1_n_0;
  wire start_count_reg_i_2_n_0;
  wire start_count_reg_i_3_n_0;
  wire start_count_reg_i_4_n_0;
  wire start_count_reg_i_5_n_0;
  wire start_count_reg_i_6_n_0;
  wire start_count_reg_i_7_n_0;
  wire start_count_reg_i_8_n_0;
  wire start_count_reg_i_9_n_0;
  wire transmit_pause_frame_valid;
  wire tx_ack0;
  wire tx_ack_reg_0;
  wire tx_ack_reg_1;
  wire tx_ack_reg_2;
  wire tx_ack_reg_3;
  wire tx_ack_reg_4;
  wire tx_ack_reg_5;
  wire tx_ack_reg_6;
  wire tx_ack_reg_7;

  (* SOFT_HLUTNM = "soft_lutpair321" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \CRC_OUT[31]_i_1__1 
       (.I0(rst_i),
        .I1(append_start_pause),
        .I2(tx_ack_reg_0),
        .O(SS));
  LUT5 #(
    .INIT(32'h0F010001)) 
    \TX_DATA_REG[10]_i_2 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [7]),
        .O(tx_ack_reg_2));
  (* SOFT_HLUTNM = "soft_lutpair315" *) 
  LUT5 #(
    .INIT(32'h0F0E000E)) 
    \TX_DATA_REG[11]_i_2 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [8]),
        .O(tx_ack_reg_4));
  LUT5 #(
    .INIT(32'h0F0E000E)) 
    \TX_DATA_REG[13]_i_2 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [9]),
        .O(tx_ack_reg_5));
  LUT5 #(
    .INIT(32'h0F0E000E)) 
    \TX_DATA_REG[15]_i_2 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [10]),
        .O(tx_ack_reg_6));
  LUT6 #(
    .INIT(64'hE2E2E2E2C0C0C0F3)) 
    \TX_DATA_REG[2]_i_1 
       (.I0(\TX_DATA_REG_reg[40] [0]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[63]_1 [0]),
        .I3(append_start_pause),
        .I4(tx_ack_reg_0),
        .I5(transmit_pause_frame_valid),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT5 #(
    .INIT(32'h0F0E000E)) 
    \TX_DATA_REG[31]_i_3 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [11]),
        .O(tx_ack_reg_7));
  LUT6 #(
    .INIT(64'hE2E2E2E2F3F3F3C0)) 
    \TX_DATA_REG[3]_i_1 
       (.I0(\TX_DATA_REG_reg[40] [1]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[63]_1 [1]),
        .I3(append_start_pause),
        .I4(tx_ack_reg_0),
        .I5(transmit_pause_frame_valid),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT5 #(
    .INIT(32'h0F010001)) 
    \TX_DATA_REG[48]_i_2 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [11]),
        .O(tx_ack_reg_3));
  LUT6 #(
    .INIT(64'hE2E2E2E2F3F3F3C0)) 
    \TX_DATA_REG[4]_i_1 
       (.I0(\TX_DATA_REG_reg[40] [2]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[63]_1 [2]),
        .I3(append_start_pause),
        .I4(tx_ack_reg_0),
        .I5(transmit_pause_frame_valid),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[58]_i_1 
       (.I0(append_start_pause_reg_0),
        .I1(\TX_DATA_REG_reg[63] ),
        .I2(\TX_DATA_REG_reg[63]_0 [0]),
        .I3(\TX_DATA_REG_reg[63]_0 [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[63]_1 [6]),
        .O(D[6]));
  (* SOFT_HLUTNM = "soft_lutpair314" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \TX_DATA_REG[58]_i_2 
       (.I0(append_start_pause),
        .I1(tx_ack_reg_0),
        .I2(transmit_pause_frame_valid),
        .I3(FRAME_START),
        .O(append_start_pause_reg_0));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[59]_i_1 
       (.I0(append_start_pause_reg),
        .I1(\TX_DATA_REG_reg[63] ),
        .I2(\TX_DATA_REG_reg[63]_0 [0]),
        .I3(\TX_DATA_REG_reg[63]_0 [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[63]_1 [7]),
        .O(D[7]));
  LUT6 #(
    .INIT(64'hE2E2E2E2F3F3F3C0)) 
    \TX_DATA_REG[5]_i_1 
       (.I0(\TX_DATA_REG_reg[40] [3]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[63]_1 [3]),
        .I3(append_start_pause),
        .I4(tx_ack_reg_0),
        .I5(transmit_pause_frame_valid),
        .O(D[3]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[61]_i_1 
       (.I0(append_start_pause_reg),
        .I1(\TX_DATA_REG_reg[63] ),
        .I2(\TX_DATA_REG_reg[63]_0 [0]),
        .I3(\TX_DATA_REG_reg[63]_0 [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[63]_1 [8]),
        .O(D[8]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[63]_i_2 
       (.I0(append_start_pause_reg),
        .I1(\TX_DATA_REG_reg[63] ),
        .I2(\TX_DATA_REG_reg[63]_0 [0]),
        .I3(\TX_DATA_REG_reg[63]_0 [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[63]_1 [9]),
        .O(D[9]));
  (* SOFT_HLUTNM = "soft_lutpair315" *) 
  LUT4 #(
    .INIT(16'h000E)) 
    \TX_DATA_REG[63]_i_5 
       (.I0(append_start_pause),
        .I1(tx_ack_reg_0),
        .I2(transmit_pause_frame_valid),
        .I3(FRAME_START),
        .O(append_start_pause_reg));
  LUT6 #(
    .INIT(64'hE2E2E2E2F3F3F3C0)) 
    \TX_DATA_REG[6]_i_1 
       (.I0(\TX_DATA_REG_reg[40] [4]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[63]_1 [4]),
        .I3(append_start_pause),
        .I4(tx_ack_reg_0),
        .I5(transmit_pause_frame_valid),
        .O(D[4]));
  LUT6 #(
    .INIT(64'hE2E2E2E2F3F3F3C0)) 
    \TX_DATA_REG[7]_i_1 
       (.I0(\TX_DATA_REG_reg[40] [5]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[63]_1 [5]),
        .I3(append_start_pause),
        .I4(tx_ack_reg_0),
        .I5(transmit_pause_frame_valid),
        .O(D[5]));
  (* SOFT_HLUTNM = "soft_lutpair314" *) 
  LUT5 #(
    .INIT(32'h0F010001)) 
    \TX_DATA_REG[8]_i_2 
       (.I0(tx_ack_reg_0),
        .I1(append_start_pause),
        .I2(FRAME_START),
        .I3(transmit_pause_frame_valid),
        .I4(\TX_DATA_REG_reg[40] [6]),
        .O(tx_ack_reg_1));
  (* SOFT_HLUTNM = "soft_lutpair322" *) 
  LUT2 #(
    .INIT(4'h2)) 
    apply_pause_delay_i_1
       (.I0(apply_pause_delay_reg),
        .I1(tx_ack_reg_0),
        .O(apply_pause_delay));
  (* SOFT_HLUTNM = "soft_lutpair316" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \counter[0]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[0]),
        .O(p_0_in[0]));
  (* SOFT_HLUTNM = "soft_lutpair319" *) 
  LUT3 #(
    .INIT(8'h82)) 
    \counter[10]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[10]_i_2_n_0 ),
        .I2(counter_reg[10]),
        .O(p_0_in[10]));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \counter[10]_i_2 
       (.I0(counter_reg[8]),
        .I1(counter_reg[6]),
        .I2(\counter[9]_i_2_n_0 ),
        .I3(counter_reg[7]),
        .I4(counter_reg[9]),
        .O(\counter[10]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair317" *) 
  LUT3 #(
    .INIT(8'h82)) 
    \counter[11]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[14]_i_2_n_0 ),
        .I2(counter_reg[11]),
        .O(p_0_in[11]));
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT4 #(
    .INIT(16'h8A20)) 
    \counter[12]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[14]_i_2_n_0 ),
        .I2(counter_reg[11]),
        .I3(counter_reg[12]),
        .O(p_0_in[12]));
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT5 #(
    .INIT(32'hA2AA0800)) 
    \counter[13]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[11]),
        .I2(\counter[14]_i_2_n_0 ),
        .I3(counter_reg[12]),
        .I4(counter_reg[13]),
        .O(p_0_in[13]));
  LUT6 #(
    .INIT(64'hAA2AAAAA00800000)) 
    \counter[14]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[13]),
        .I2(counter_reg[12]),
        .I3(\counter[14]_i_2_n_0 ),
        .I4(counter_reg[11]),
        .I5(counter_reg[14]),
        .O(p_0_in[14]));
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \counter[14]_i_2 
       (.I0(counter_reg[9]),
        .I1(counter_reg[7]),
        .I2(\counter[9]_i_2_n_0 ),
        .I3(counter_reg[6]),
        .I4(counter_reg[8]),
        .I5(counter_reg[10]),
        .O(\counter[14]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \counter[15]_i_1__0 
       (.I0(start_count),
        .I1(start_count_reg_i_3_n_0),
        .O(\counter[15]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair316" *) 
  LUT4 #(
    .INIT(16'h2A80)) 
    \counter[15]_i_2 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[15]_i_3_n_0 ),
        .I2(counter_reg[14]),
        .I3(counter_reg[15]),
        .O(p_0_in[15]));
  (* SOFT_HLUTNM = "soft_lutpair320" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \counter[15]_i_2__0 
       (.I0(tx_ack_reg_0),
        .I1(rst_i),
        .O(AR));
  (* SOFT_HLUTNM = "soft_lutpair317" *) 
  LUT4 #(
    .INIT(16'h0800)) 
    \counter[15]_i_3 
       (.I0(counter_reg[13]),
        .I1(counter_reg[12]),
        .I2(\counter[14]_i_2_n_0 ),
        .I3(counter_reg[11]),
        .O(\counter[15]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair318" *) 
  LUT3 #(
    .INIT(8'h28)) 
    \counter[1]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[0]),
        .I2(counter_reg[1]),
        .O(p_0_in[1]));
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT4 #(
    .INIT(16'h2A80)) 
    \counter[2]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[1]),
        .I2(counter_reg[0]),
        .I3(counter_reg[2]),
        .O(p_0_in[2]));
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    \counter[3]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[0]),
        .I2(counter_reg[1]),
        .I3(counter_reg[2]),
        .I4(counter_reg[3]),
        .O(p_0_in[3]));
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    \counter[4]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[2]),
        .I2(counter_reg[1]),
        .I3(counter_reg[0]),
        .I4(counter_reg[3]),
        .I5(counter_reg[4]),
        .O(p_0_in[4]));
  (* SOFT_HLUTNM = "soft_lutpair318" *) 
  LUT3 #(
    .INIT(8'h82)) 
    \counter[5]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[5]_i_2_n_0 ),
        .I2(counter_reg[5]),
        .O(p_0_in[5]));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \counter[5]_i_2 
       (.I0(counter_reg[3]),
        .I1(counter_reg[0]),
        .I2(counter_reg[1]),
        .I3(counter_reg[2]),
        .I4(counter_reg[4]),
        .O(\counter[5]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair319" *) 
  LUT3 #(
    .INIT(8'h82)) 
    \counter[6]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[9]_i_2_n_0 ),
        .I2(counter_reg[6]),
        .O(p_0_in[6]));
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT4 #(
    .INIT(16'h8A20)) 
    \counter[7]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(\counter[9]_i_2_n_0 ),
        .I2(counter_reg[6]),
        .I3(counter_reg[7]),
        .O(p_0_in[7]));
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT5 #(
    .INIT(32'hA2AA0800)) 
    \counter[8]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[6]),
        .I2(\counter[9]_i_2_n_0 ),
        .I3(counter_reg[7]),
        .I4(counter_reg[8]),
        .O(p_0_in[8]));
  LUT6 #(
    .INIT(64'hA2AAAAAA08000000)) 
    \counter[9]_i_1__0 
       (.I0(start_count_reg_i_3_n_0),
        .I1(counter_reg[7]),
        .I2(\counter[9]_i_2_n_0 ),
        .I3(counter_reg[6]),
        .I4(counter_reg[8]),
        .I5(counter_reg[9]),
        .O(p_0_in[9]));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \counter[9]_i_2 
       (.I0(counter_reg[4]),
        .I1(counter_reg[2]),
        .I2(counter_reg[1]),
        .I3(counter_reg[0]),
        .I4(counter_reg[3]),
        .I5(counter_reg[5]),
        .O(\counter[9]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[0] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[0]),
        .Q(counter_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[10] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[10]),
        .Q(counter_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[11] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[11]),
        .Q(counter_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[12] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[12]),
        .Q(counter_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[13] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[13]),
        .Q(counter_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[14] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[14]),
        .Q(counter_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[15] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[15]),
        .Q(counter_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[1] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[1]),
        .Q(counter_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[2] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[2]),
        .Q(counter_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[3] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[3]),
        .Q(counter_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[4] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[4]),
        .Q(counter_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[5] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[5]),
        .Q(counter_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[6] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[6]),
        .Q(counter_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[7] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[7]),
        .Q(counter_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[8] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[8]),
        .Q(counter_reg[8]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[9] 
       (.C(clk_i),
        .CE(\counter[15]_i_1__0_n_0 ),
        .CLR(reset0),
        .D(p_0_in[9]),
        .Q(counter_reg[9]));
  LUT2 #(
    .INIT(4'hE)) 
    start_count_del_i_1
       (.I0(reset_tx_int),
        .I1(rst_i),
        .O(reset0));
  FDCE #(
    .INIT(1'b0)) 
    start_count_del_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset0),
        .D(start_count),
        .Q(start_count_del));
  LDCE #(
    .INIT(1'b0)) 
    start_count_reg
       (.CLR(1'b0),
        .D(start_count_reg_i_1_n_0),
        .G(start_count_reg_i_2_n_0),
        .GE(1'b1),
        .Q(start_count));
  (* SOFT_HLUTNM = "soft_lutpair320" *) 
  LUT3 #(
    .INIT(8'h02)) 
    start_count_reg_i_1
       (.I0(out),
        .I1(rst_i),
        .I2(reset_tx_int),
        .O(start_count_reg_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEEEF)) 
    start_count_reg_i_2
       (.I0(reset_tx_int),
        .I1(rst_i),
        .I2(start_count_reg_i_3_n_0),
        .I3(FRAME_START),
        .I4(start_count_del_reg_0),
        .I5(out),
        .O(start_count_reg_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    start_count_reg_i_3
       (.I0(start_count_reg_i_4_n_0),
        .I1(start_count_reg_i_5_n_0),
        .I2(start_count_reg_i_6_n_0),
        .I3(start_count_reg_i_7_n_0),
        .I4(start_count_reg_i_8_n_0),
        .I5(start_count_reg_i_9_n_0),
        .O(start_count_reg_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    start_count_reg_i_4
       (.I0(Q[14]),
        .I1(counter_reg[14]),
        .I2(counter_reg[13]),
        .I3(Q[13]),
        .I4(counter_reg[12]),
        .I5(Q[12]),
        .O(start_count_reg_i_4_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    start_count_reg_i_5
       (.I0(Q[6]),
        .I1(counter_reg[6]),
        .I2(counter_reg[7]),
        .I3(Q[7]),
        .I4(counter_reg[8]),
        .I5(Q[8]),
        .O(start_count_reg_i_5_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    start_count_reg_i_6
       (.I0(Q[9]),
        .I1(counter_reg[9]),
        .I2(counter_reg[11]),
        .I3(Q[11]),
        .I4(counter_reg[10]),
        .I5(Q[10]),
        .O(start_count_reg_i_6_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    start_count_reg_i_7
       (.I0(Q[3]),
        .I1(counter_reg[3]),
        .I2(counter_reg[4]),
        .I3(Q[4]),
        .I4(counter_reg[5]),
        .I5(Q[5]),
        .O(start_count_reg_i_7_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    start_count_reg_i_8
       (.I0(Q[2]),
        .I1(counter_reg[2]),
        .I2(counter_reg[1]),
        .I3(Q[1]),
        .I4(counter_reg[0]),
        .I5(Q[0]),
        .O(start_count_reg_i_8_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    start_count_reg_i_9
       (.I0(counter_reg[15]),
        .I1(Q[15]),
        .O(start_count_reg_i_9_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[0]_i_1 
       (.I0(I94[0]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [0]));
  (* SOFT_HLUTNM = "soft_lutpair325" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[10]_i_1 
       (.I0(I94[10]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [10]));
  (* SOFT_HLUTNM = "soft_lutpair324" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[11]_i_1 
       (.I0(I94[11]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [11]));
  (* SOFT_HLUTNM = "soft_lutpair324" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[12]_i_1 
       (.I0(I94[12]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [12]));
  (* SOFT_HLUTNM = "soft_lutpair323" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[13]_i_1 
       (.I0(I94[13]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [13]));
  (* SOFT_HLUTNM = "soft_lutpair323" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[14]_i_1 
       (.I0(I94[14]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [14]));
  (* SOFT_HLUTNM = "soft_lutpair321" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \store_pause_frame[15]_i_1 
       (.I0(tx_ack_reg_0),
        .I1(apply_pause_delay_reg),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair322" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[15]_i_2 
       (.I0(I94[15]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [15]));
  (* SOFT_HLUTNM = "soft_lutpair329" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[1]_i_1 
       (.I0(I94[1]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [1]));
  (* SOFT_HLUTNM = "soft_lutpair329" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[2]_i_1 
       (.I0(I94[2]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [2]));
  (* SOFT_HLUTNM = "soft_lutpair328" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[3]_i_1 
       (.I0(I94[3]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [3]));
  (* SOFT_HLUTNM = "soft_lutpair328" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[4]_i_1 
       (.I0(I94[4]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [4]));
  (* SOFT_HLUTNM = "soft_lutpair327" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[5]_i_1 
       (.I0(I94[5]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [5]));
  (* SOFT_HLUTNM = "soft_lutpair327" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[6]_i_1 
       (.I0(I94[6]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [6]));
  (* SOFT_HLUTNM = "soft_lutpair326" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[7]_i_1 
       (.I0(I94[7]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [7]));
  (* SOFT_HLUTNM = "soft_lutpair326" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[8]_i_1 
       (.I0(I94[8]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [8]));
  (* SOFT_HLUTNM = "soft_lutpair325" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \store_pause_frame[9]_i_1 
       (.I0(I94[9]),
        .I1(tx_ack_reg_0),
        .O(\FC_TX_PAUSEDATA_reg[15] [9]));
  LUT2 #(
    .INIT(4'h2)) 
    tx_ack_i_1
       (.I0(start_count_del),
        .I1(start_count),
        .O(tx_ack0));
  FDCE #(
    .INIT(1'b0)) 
    tx_ack_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset0),
        .D(tx_ack0),
        .Q(tx_ack_reg_0));
endmodule

(* ORIG_REF_NAME = "byte_count_module" *) 
module switch_elements_byte_count_module
   (Q,
    D,
    \TX_DATA_REG_reg[15] ,
    E,
    \enable_i[6] ,
    \TX_DATA_VALID_DELAY_reg[62] ,
    \BYTE_COUNTER_reg[3]_0 ,
    \BYTE_COUNTER_reg[3]_1 ,
    tx_ack_reg,
    vlan_enabled_int,
    \final_byte_count_reg[15] ,
    load_CRC8,
    \final_byte_count_reg[15]_0 ,
    \final_byte_count_reg[3] ,
    \final_byte_count_reg[4] ,
    \final_byte_count_reg[5] ,
    \final_byte_count_reg[6] ,
    \final_byte_count_reg[8] ,
    \final_byte_count_reg[9] ,
    \final_byte_count_reg[10] ,
    \final_byte_count_reg[11] ,
    \final_byte_count_reg[13] ,
    \final_byte_count_reg[14] ,
    \length_register_reg[15] ,
    out,
    \TX_DATA_VALID_REG_reg[7] ,
    FRAME_START,
    transmit_pause_frame_del,
    \TX_DATA_VALID_REG_reg[4] ,
    \TX_DATA_REG_reg[16] ,
    \TX_DATA_REG_reg[62] ,
    \TX_DATA_REG_reg[62]_0 ,
    transmit_pause_frame_valid,
    \TX_DATA_REG_reg[19] ,
    \TX_DATA_REG_reg[20] ,
    \TX_DATA_REG_reg[21] ,
    \TX_DATA_REG_reg[33] ,
    \TX_DATA_REG_reg[40] ,
    \TX_DATA_REG_reg[15]_0 ,
    \TX_DATA_REG_reg[14] ,
    \TX_DATA_REG_reg[13] ,
    \TX_DATA_REG_reg[12] ,
    \TX_DATA_REG_reg[11] ,
    \TX_DATA_REG_reg[10] ,
    \TX_DATA_REG_reg[9] ,
    \TX_DATA_REG_reg[8] ,
    \TX_DATA_REG_reg[0] ,
    frame_start_del,
    TX_ACK,
    FRAME_START_reg,
    clk_i,
    AR);
  output [13:0]Q;
  output [13:0]D;
  output [15:0]\TX_DATA_REG_reg[15] ;
  output [0:0]E;
  output [7:0]\enable_i[6] ;
  output [51:0]\TX_DATA_VALID_DELAY_reg[62] ;
  output \BYTE_COUNTER_reg[3]_0 ;
  output [0:0]\BYTE_COUNTER_reg[3]_1 ;
  output tx_ack_reg;
  input vlan_enabled_int;
  input [13:0]\final_byte_count_reg[15] ;
  input load_CRC8;
  input [15:0]\final_byte_count_reg[15]_0 ;
  input \final_byte_count_reg[3] ;
  input \final_byte_count_reg[4] ;
  input \final_byte_count_reg[5] ;
  input \final_byte_count_reg[6] ;
  input \final_byte_count_reg[8] ;
  input \final_byte_count_reg[9] ;
  input \final_byte_count_reg[10] ;
  input \final_byte_count_reg[11] ;
  input \final_byte_count_reg[13] ;
  input \final_byte_count_reg[14] ;
  input [31:0]\length_register_reg[15] ;
  input out;
  input [7:0]\TX_DATA_VALID_REG_reg[7] ;
  input FRAME_START;
  input transmit_pause_frame_del;
  input [1:0]\TX_DATA_VALID_REG_reg[4] ;
  input \TX_DATA_REG_reg[16] ;
  input [7:0]\TX_DATA_REG_reg[62] ;
  input [51:0]\TX_DATA_REG_reg[62]_0 ;
  input transmit_pause_frame_valid;
  input \TX_DATA_REG_reg[19] ;
  input \TX_DATA_REG_reg[20] ;
  input \TX_DATA_REG_reg[21] ;
  input \TX_DATA_REG_reg[33] ;
  input \TX_DATA_REG_reg[40] ;
  input \TX_DATA_REG_reg[15]_0 ;
  input \TX_DATA_REG_reg[14] ;
  input \TX_DATA_REG_reg[13] ;
  input \TX_DATA_REG_reg[12] ;
  input \TX_DATA_REG_reg[11] ;
  input \TX_DATA_REG_reg[10] ;
  input \TX_DATA_REG_reg[9] ;
  input \TX_DATA_REG_reg[8] ;
  input \TX_DATA_REG_reg[0] ;
  input frame_start_del;
  input TX_ACK;
  input FRAME_START_reg;
  input clk_i;
  input [0:0]AR;

  wire [0:0]AR;
  wire \BYTE_COUNTER_reg[3]_0 ;
  wire [0:0]\BYTE_COUNTER_reg[3]_1 ;
  wire [13:0]D;
  wire [0:0]E;
  wire FRAME_START;
  wire FRAME_START_i_2_n_0;
  wire FRAME_START_reg;
  wire [13:0]Q;
  wire START0;
  wire TX_ACK;
  wire \TX_DATA_REG[23]_i_2_n_0 ;
  wire \TX_DATA_REG[31]_i_2_n_0 ;
  wire \TX_DATA_REG[39]_i_2_n_0 ;
  wire \TX_DATA_REG[47]_i_2_n_0 ;
  wire \TX_DATA_REG[55]_i_2_n_0 ;
  wire \TX_DATA_REG[55]_i_3_n_0 ;
  wire \TX_DATA_REG[55]_i_4_n_0 ;
  wire \TX_DATA_REG[55]_i_5_n_0 ;
  wire \TX_DATA_REG_reg[0] ;
  wire \TX_DATA_REG_reg[10] ;
  wire \TX_DATA_REG_reg[11] ;
  wire \TX_DATA_REG_reg[12] ;
  wire \TX_DATA_REG_reg[13] ;
  wire \TX_DATA_REG_reg[14] ;
  wire [15:0]\TX_DATA_REG_reg[15] ;
  wire \TX_DATA_REG_reg[15]_0 ;
  wire \TX_DATA_REG_reg[16] ;
  wire \TX_DATA_REG_reg[19] ;
  wire \TX_DATA_REG_reg[20] ;
  wire \TX_DATA_REG_reg[21] ;
  wire \TX_DATA_REG_reg[33] ;
  wire \TX_DATA_REG_reg[40] ;
  wire [7:0]\TX_DATA_REG_reg[62] ;
  wire [51:0]\TX_DATA_REG_reg[62]_0 ;
  wire \TX_DATA_REG_reg[8] ;
  wire \TX_DATA_REG_reg[9] ;
  wire [51:0]\TX_DATA_VALID_DELAY_reg[62] ;
  wire \TX_DATA_VALID_REG[3]_i_2_n_0 ;
  wire \TX_DATA_VALID_REG[3]_i_3_n_0 ;
  wire \TX_DATA_VALID_REG[7]_i_2_n_0 ;
  wire \TX_DATA_VALID_REG[7]_i_3_n_0 ;
  wire [1:0]\TX_DATA_VALID_REG_reg[4] ;
  wire [7:0]\TX_DATA_VALID_REG_reg[7] ;
  wire clk_i;
  wire counter0_carry__0_n_3;
  wire counter0_carry__0_n_4;
  wire counter0_carry__0_n_5;
  wire counter0_carry__0_n_6;
  wire counter0_carry__0_n_7;
  wire counter0_carry_i_1_n_0;
  wire counter0_carry_n_0;
  wire counter0_carry_n_1;
  wire counter0_carry_n_2;
  wire counter0_carry_n_3;
  wire counter0_carry_n_4;
  wire counter0_carry_n_5;
  wire counter0_carry_n_6;
  wire counter0_carry_n_7;
  wire [15:2]counter_reg;
  wire [7:0]\enable_i[6] ;
  wire \final_byte_count[15]_i_2_n_0 ;
  wire \final_byte_count[15]_i_4_n_0 ;
  wire \final_byte_count[15]_i_5_n_0 ;
  wire \final_byte_count[5]_i_2_n_0 ;
  wire \final_byte_count[5]_i_4_n_0 ;
  wire \final_byte_count_reg[10] ;
  wire \final_byte_count_reg[11] ;
  wire \final_byte_count_reg[13] ;
  wire \final_byte_count_reg[14] ;
  wire [13:0]\final_byte_count_reg[15] ;
  wire [15:0]\final_byte_count_reg[15]_0 ;
  wire \final_byte_count_reg[3] ;
  wire \final_byte_count_reg[4] ;
  wire \final_byte_count_reg[5] ;
  wire \final_byte_count_reg[6] ;
  wire \final_byte_count_reg[8] ;
  wire \final_byte_count_reg[9] ;
  wire frame_start_del;
  wire \length_register[15]_i_3_n_0 ;
  wire \length_register[15]_i_4_n_0 ;
  wire \length_register[15]_i_5_n_0 ;
  wire [31:0]\length_register_reg[15] ;
  wire load_CRC8;
  wire out;
  wire [15:2]p_0_in__1;
  wire transmit_pause_frame_del;
  wire transmit_pause_frame_valid;
  wire tx_ack_reg;
  wire vlan_enabled_int;
  wire [7:5]NLW_counter0_carry__0_CO_UNCONNECTED;
  wire [7:6]NLW_counter0_carry__0_O_UNCONNECTED;

  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[10]),
        .Q(Q[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[11]),
        .Q(Q[9]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[12]),
        .Q(Q[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[13]),
        .Q(Q[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[14]),
        .Q(Q[12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[15]),
        .Q(Q[13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[2]),
        .Q(Q[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[3]),
        .Q(Q[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[4]),
        .Q(Q[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[5]),
        .Q(Q[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[6]),
        .Q(Q[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[7]),
        .Q(Q[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[8]),
        .Q(Q[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \BYTE_COUNTER_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(counter_reg[9]),
        .Q(Q[7]),
        .R(1'b0));
  LUT6 #(
    .INIT(64'hABAAFFFFAAAAAAAA)) 
    FRAME_START_i_1
       (.I0(TX_ACK),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(FRAME_START_i_2_n_0),
        .I4(FRAME_START_reg),
        .I5(FRAME_START),
        .O(tx_ack_reg));
  (* SOFT_HLUTNM = "soft_lutpair408" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    FRAME_START_i_2
       (.I0(Q[4]),
        .I1(Q[5]),
        .I2(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I3(Q[1]),
        .I4(Q[0]),
        .O(FRAME_START_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[10]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [2]),
        .I5(\TX_DATA_REG_reg[10] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[11]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [3]),
        .I5(\TX_DATA_REG_reg[11] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [3]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[12]_i_1 
       (.I0(\TX_DATA_REG_reg[12] ),
        .I1(\BYTE_COUNTER_reg[3]_0 ),
        .I2(\TX_DATA_REG_reg[62] [0]),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[62]_0 [4]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[13]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [5]),
        .I5(\TX_DATA_REG_reg[13] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [5]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[14]_i_1 
       (.I0(\TX_DATA_REG_reg[14] ),
        .I1(\BYTE_COUNTER_reg[3]_0 ),
        .I2(\TX_DATA_REG_reg[62] [0]),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[62]_0 [6]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[15]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [7]),
        .I5(\TX_DATA_REG_reg[15]_0 ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [7]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[16]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[23]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [8]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [8]));
  LUT6 #(
    .INIT(64'h05050505C5C5C505)) 
    \TX_DATA_REG[17]_i_1 
       (.I0(transmit_pause_frame_valid),
        .I1(\TX_DATA_REG_reg[62]_0 [9]),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG[23]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [9]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[18]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[23]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [10]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [10]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[19]_i_1 
       (.I0(\TX_DATA_REG_reg[19] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[23]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [11]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [11]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[20]_i_1 
       (.I0(\TX_DATA_REG_reg[20] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[23]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [12]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [12]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[21]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[23]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [13]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [13]));
  LUT6 #(
    .INIT(64'hAA80AA8A00000000)) 
    \TX_DATA_REG[22]_i_1 
       (.I0(\TX_DATA_REG_reg[62]_0 [14]),
        .I1(\TX_DATA_REG_reg[62] [2]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\BYTE_COUNTER_reg[3]_0 ),
        .I4(\TX_DATA_REG_reg[62] [0]),
        .I5(FRAME_START),
        .O(\TX_DATA_VALID_DELAY_reg[62] [14]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[23]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[23]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [15]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [15]));
  LUT6 #(
    .INIT(64'h0000040004000400)) 
    \TX_DATA_REG[23]_i_2 
       (.I0(\TX_DATA_REG_reg[62] [2]),
        .I1(\TX_DATA_REG_reg[62] [1]),
        .I2(\TX_DATA_REG[55]_i_4_n_0 ),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(\TX_DATA_REG[55]_i_5_n_0 ),
        .I5(Q[1]),
        .O(\TX_DATA_REG[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[24]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[31]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [16]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [16]));
  LUT6 #(
    .INIT(64'h05050505C5C5C505)) 
    \TX_DATA_REG[25]_i_1 
       (.I0(transmit_pause_frame_valid),
        .I1(\TX_DATA_REG_reg[62]_0 [17]),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG[31]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [17]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[26]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[31]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [18]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [18]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[27]_i_1 
       (.I0(\TX_DATA_REG_reg[19] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[31]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [19]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [19]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[28]_i_1 
       (.I0(\TX_DATA_REG_reg[20] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[31]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [20]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [20]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[29]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[31]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [21]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [21]));
  LUT6 #(
    .INIT(64'hAA80AA8A00000000)) 
    \TX_DATA_REG[30]_i_1 
       (.I0(\TX_DATA_REG_reg[62]_0 [22]),
        .I1(\TX_DATA_REG_reg[62] [3]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\BYTE_COUNTER_reg[3]_0 ),
        .I4(\TX_DATA_REG_reg[62] [0]),
        .I5(FRAME_START),
        .O(\TX_DATA_VALID_DELAY_reg[62] [22]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00A80000)) 
    \TX_DATA_REG[31]_i_1 
       (.I0(FRAME_START),
        .I1(\TX_DATA_REG_reg[62] [1]),
        .I2(\TX_DATA_REG[55]_i_3_n_0 ),
        .I3(\TX_DATA_REG[31]_i_2_n_0 ),
        .I4(\TX_DATA_REG_reg[62]_0 [23]),
        .I5(\TX_DATA_REG_reg[19] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [23]));
  LUT6 #(
    .INIT(64'h0000040004000400)) 
    \TX_DATA_REG[31]_i_2 
       (.I0(\TX_DATA_REG_reg[62] [3]),
        .I1(\TX_DATA_REG_reg[62] [1]),
        .I2(\TX_DATA_REG[55]_i_4_n_0 ),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(\TX_DATA_REG[55]_i_5_n_0 ),
        .I5(Q[1]),
        .O(\TX_DATA_REG[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[32]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [24]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [24]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[33]_i_1 
       (.I0(\TX_DATA_REG_reg[33] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [25]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [25]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[34]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [26]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [26]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[35]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [27]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [27]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[36]_i_1 
       (.I0(\TX_DATA_REG_reg[20] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [28]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [28]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[37]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [29]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [29]));
  LUT6 #(
    .INIT(64'hAA80AA8A00000000)) 
    \TX_DATA_REG[38]_i_1 
       (.I0(\TX_DATA_REG_reg[62]_0 [30]),
        .I1(\TX_DATA_REG_reg[62] [4]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\BYTE_COUNTER_reg[3]_0 ),
        .I4(\TX_DATA_REG_reg[62] [0]),
        .I5(FRAME_START),
        .O(\TX_DATA_VALID_DELAY_reg[62] [30]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[39]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[39]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [31]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [31]));
  LUT6 #(
    .INIT(64'h0000040004000400)) 
    \TX_DATA_REG[39]_i_2 
       (.I0(\TX_DATA_REG_reg[62] [4]),
        .I1(\TX_DATA_REG_reg[62] [1]),
        .I2(\TX_DATA_REG[55]_i_4_n_0 ),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(\TX_DATA_REG[55]_i_5_n_0 ),
        .I5(Q[1]),
        .O(\TX_DATA_REG[39]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[40]_i_1 
       (.I0(\TX_DATA_REG_reg[40] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[47]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [32]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [32]));
  LUT6 #(
    .INIT(64'h05050505C5C5C505)) 
    \TX_DATA_REG[41]_i_1 
       (.I0(transmit_pause_frame_valid),
        .I1(\TX_DATA_REG_reg[62]_0 [33]),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG[47]_i_2_n_0 ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [33]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[42]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[47]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [34]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [34]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[43]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[47]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [35]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [35]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[44]_i_1 
       (.I0(\TX_DATA_REG_reg[20] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[47]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [36]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [36]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[45]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[47]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [37]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [37]));
  LUT6 #(
    .INIT(64'hAA80AA8A00000000)) 
    \TX_DATA_REG[46]_i_1 
       (.I0(\TX_DATA_REG_reg[62]_0 [38]),
        .I1(\TX_DATA_REG_reg[62] [5]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\BYTE_COUNTER_reg[3]_0 ),
        .I4(\TX_DATA_REG_reg[62] [0]),
        .I5(FRAME_START),
        .O(\TX_DATA_VALID_DELAY_reg[62] [38]));
  LUT6 #(
    .INIT(64'hAAAAEEEAAAAAAAAA)) 
    \TX_DATA_REG[47]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG[47]_i_2_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [39]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [39]));
  LUT6 #(
    .INIT(64'h0000040004000400)) 
    \TX_DATA_REG[47]_i_2 
       (.I0(\TX_DATA_REG_reg[62] [5]),
        .I1(\TX_DATA_REG_reg[62] [1]),
        .I2(\TX_DATA_REG[55]_i_4_n_0 ),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(\TX_DATA_REG[55]_i_5_n_0 ),
        .I5(Q[1]),
        .O(\TX_DATA_REG[47]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF44400000)) 
    \TX_DATA_REG[48]_i_1 
       (.I0(\TX_DATA_REG[55]_i_2_n_0 ),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(\TX_DATA_REG[55]_i_3_n_0 ),
        .I4(\TX_DATA_REG_reg[62]_0 [40]),
        .I5(\TX_DATA_REG_reg[40] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [40]));
  LUT6 #(
    .INIT(64'h0C550C550C550055)) 
    \TX_DATA_REG[49]_i_1 
       (.I0(transmit_pause_frame_valid),
        .I1(\TX_DATA_REG_reg[62]_0 [41]),
        .I2(\TX_DATA_REG[55]_i_2_n_0 ),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62] [1]),
        .I5(\TX_DATA_REG[55]_i_3_n_0 ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [41]));
  LUT6 #(
    .INIT(64'hBABABAAAAAAAAAAA)) 
    \TX_DATA_REG[50]_i_1 
       (.I0(\TX_DATA_REG_reg[16] ),
        .I1(\TX_DATA_REG[55]_i_2_n_0 ),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [42]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [42]));
  LUT6 #(
    .INIT(64'hBABABAAAAAAAAAAA)) 
    \TX_DATA_REG[51]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(\TX_DATA_REG[55]_i_2_n_0 ),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [43]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [43]));
  LUT6 #(
    .INIT(64'hBABABAAAAAAAAAAA)) 
    \TX_DATA_REG[52]_i_1 
       (.I0(\TX_DATA_REG_reg[20] ),
        .I1(\TX_DATA_REG[55]_i_2_n_0 ),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [44]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [44]));
  LUT6 #(
    .INIT(64'hBABABAAAAAAAAAAA)) 
    \TX_DATA_REG[53]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(\TX_DATA_REG[55]_i_2_n_0 ),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [45]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [45]));
  LUT6 #(
    .INIT(64'hAA8A0000888A0000)) 
    \TX_DATA_REG[54]_i_1 
       (.I0(\TX_DATA_REG_reg[62]_0 [46]),
        .I1(\BYTE_COUNTER_reg[3]_0 ),
        .I2(\TX_DATA_REG_reg[62] [0]),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[62] [6]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [46]));
  LUT6 #(
    .INIT(64'hBABABAAAAAAAAAAA)) 
    \TX_DATA_REG[55]_i_1 
       (.I0(\TX_DATA_REG_reg[21] ),
        .I1(\TX_DATA_REG[55]_i_2_n_0 ),
        .I2(FRAME_START),
        .I3(\TX_DATA_REG_reg[62] [1]),
        .I4(\TX_DATA_REG[55]_i_3_n_0 ),
        .I5(\TX_DATA_REG_reg[62]_0 [47]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [47]));
  LUT6 #(
    .INIT(64'h0000040004000400)) 
    \TX_DATA_REG[55]_i_2 
       (.I0(\TX_DATA_REG_reg[62] [6]),
        .I1(\TX_DATA_REG_reg[62] [1]),
        .I2(\TX_DATA_REG[55]_i_4_n_0 ),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(\TX_DATA_REG[55]_i_5_n_0 ),
        .I5(Q[1]),
        .O(\TX_DATA_REG[55]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFBBBBBBBFFFFFFFF)) 
    \TX_DATA_REG[55]_i_3 
       (.I0(\TX_DATA_REG[55]_i_4_n_0 ),
        .I1(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I2(Q[3]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(\TX_DATA_REG_reg[62] [0]),
        .O(\TX_DATA_REG[55]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair409" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \TX_DATA_REG[55]_i_4 
       (.I0(Q[4]),
        .I1(Q[5]),
        .O(\TX_DATA_REG[55]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \TX_DATA_REG[55]_i_5 
       (.I0(Q[2]),
        .I1(Q[3]),
        .O(\TX_DATA_REG[55]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[56]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [7]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [48]),
        .I5(\TX_DATA_REG_reg[33] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [48]));
  LUT6 #(
    .INIT(64'hCCCCC0CC55555555)) 
    \TX_DATA_REG[57]_i_1 
       (.I0(transmit_pause_frame_valid),
        .I1(\TX_DATA_REG_reg[62]_0 [49]),
        .I2(\BYTE_COUNTER_reg[3]_0 ),
        .I3(\TX_DATA_REG_reg[62] [0]),
        .I4(\TX_DATA_REG_reg[62] [7]),
        .I5(FRAME_START),
        .O(\TX_DATA_VALID_DELAY_reg[62] [49]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \TX_DATA_REG[60]_i_1 
       (.I0(\TX_DATA_REG_reg[20] ),
        .I1(\BYTE_COUNTER_reg[3]_0 ),
        .I2(\TX_DATA_REG_reg[62] [0]),
        .I3(\TX_DATA_REG_reg[62] [7]),
        .I4(FRAME_START),
        .I5(\TX_DATA_REG_reg[62]_0 [50]),
        .O(\TX_DATA_VALID_DELAY_reg[62] [50]));
  LUT5 #(
    .INIT(32'h88888088)) 
    \TX_DATA_REG[62]_i_1 
       (.I0(\TX_DATA_REG_reg[62]_0 [51]),
        .I1(FRAME_START),
        .I2(\TX_DATA_REG_reg[62] [7]),
        .I3(\TX_DATA_REG_reg[62] [0]),
        .I4(\BYTE_COUNTER_reg[3]_0 ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [51]));
  LUT2 #(
    .INIT(4'hE)) 
    \TX_DATA_REG[63]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[0] ),
        .O(\BYTE_COUNTER_reg[3]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF80FF)) 
    \TX_DATA_REG[63]_i_3 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(Q[5]),
        .I5(Q[4]),
        .O(\BYTE_COUNTER_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[8]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [0]),
        .I5(\TX_DATA_REG_reg[8] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \TX_DATA_REG[9]_i_1 
       (.I0(\BYTE_COUNTER_reg[3]_0 ),
        .I1(\TX_DATA_REG_reg[62] [0]),
        .I2(\TX_DATA_REG_reg[62] [1]),
        .I3(FRAME_START),
        .I4(\TX_DATA_REG_reg[62]_0 [1]),
        .I5(\TX_DATA_REG_reg[9] ),
        .O(\TX_DATA_VALID_DELAY_reg[62] [1]));
  LUT6 #(
    .INIT(64'hBAFFBA00BA00BA00)) 
    \TX_DATA_VALID_REG[0]_i_1 
       (.I0(\TX_DATA_VALID_REG[3]_i_2_n_0 ),
        .I1(out),
        .I2(\TX_DATA_VALID_REG_reg[7] [0]),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [0]),
        .O(\enable_i[6] [0]));
  LUT6 #(
    .INIT(64'hBAFFBA00BA00BA00)) 
    \TX_DATA_VALID_REG[1]_i_1 
       (.I0(\TX_DATA_VALID_REG[3]_i_2_n_0 ),
        .I1(out),
        .I2(\TX_DATA_VALID_REG_reg[7] [1]),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [0]),
        .O(\enable_i[6] [1]));
  LUT6 #(
    .INIT(64'hBAFFBA00BA00BA00)) 
    \TX_DATA_VALID_REG[2]_i_1 
       (.I0(\TX_DATA_VALID_REG[3]_i_2_n_0 ),
        .I1(out),
        .I2(\TX_DATA_VALID_REG_reg[7] [2]),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [0]),
        .O(\enable_i[6] [2]));
  LUT6 #(
    .INIT(64'hF4FFF400F400F400)) 
    \TX_DATA_VALID_REG[3]_i_1 
       (.I0(out),
        .I1(\TX_DATA_VALID_REG_reg[7] [3]),
        .I2(\TX_DATA_VALID_REG[3]_i_2_n_0 ),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [0]),
        .O(\enable_i[6] [3]));
  LUT6 #(
    .INIT(64'h000000000000BF00)) 
    \TX_DATA_VALID_REG[3]_i_2 
       (.I0(\TX_DATA_VALID_REG[3]_i_3_n_0 ),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I4(Q[5]),
        .I5(Q[4]),
        .O(\TX_DATA_VALID_REG[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \TX_DATA_VALID_REG[3]_i_3 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\TX_DATA_VALID_REG[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBAFFBA00BA00BA00)) 
    \TX_DATA_VALID_REG[4]_i_1 
       (.I0(\TX_DATA_VALID_REG[7]_i_2_n_0 ),
        .I1(out),
        .I2(\TX_DATA_VALID_REG_reg[7] [4]),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [1]),
        .O(\enable_i[6] [4]));
  LUT6 #(
    .INIT(64'hBAFFBA00BA00BA00)) 
    \TX_DATA_VALID_REG[5]_i_1 
       (.I0(\TX_DATA_VALID_REG[7]_i_2_n_0 ),
        .I1(out),
        .I2(\TX_DATA_VALID_REG_reg[7] [5]),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [1]),
        .O(\enable_i[6] [5]));
  LUT6 #(
    .INIT(64'hBAFFBA00BA00BA00)) 
    \TX_DATA_VALID_REG[6]_i_1 
       (.I0(\TX_DATA_VALID_REG[7]_i_2_n_0 ),
        .I1(out),
        .I2(\TX_DATA_VALID_REG_reg[7] [6]),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [1]),
        .O(\enable_i[6] [6]));
  LUT6 #(
    .INIT(64'hF4FFF400F400F400)) 
    \TX_DATA_VALID_REG[7]_i_1 
       (.I0(out),
        .I1(\TX_DATA_VALID_REG_reg[7] [7]),
        .I2(\TX_DATA_VALID_REG[7]_i_2_n_0 ),
        .I3(FRAME_START),
        .I4(transmit_pause_frame_del),
        .I5(\TX_DATA_VALID_REG_reg[4] [1]),
        .O(\enable_i[6] [7]));
  (* SOFT_HLUTNM = "soft_lutpair409" *) 
  LUT5 #(
    .INIT(32'h00101010)) 
    \TX_DATA_VALID_REG[7]_i_2 
       (.I0(Q[4]),
        .I1(Q[5]),
        .I2(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I3(Q[3]),
        .I4(Q[2]),
        .O(\TX_DATA_VALID_REG[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \TX_DATA_VALID_REG[7]_i_3 
       (.I0(\final_byte_count[15]_i_5_n_0 ),
        .I1(Q[13]),
        .I2(Q[12]),
        .I3(Q[10]),
        .I4(Q[11]),
        .O(\TX_DATA_VALID_REG[7]_i_3_n_0 ));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    counter0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({counter0_carry_n_0,counter0_carry_n_1,counter0_carry_n_2,counter0_carry_n_3,counter0_carry_n_4,counter0_carry_n_5,counter0_carry_n_6,counter0_carry_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,counter_reg[3],1'b0}),
        .O(p_0_in__1[9:2]),
        .S({counter_reg[9:4],counter0_carry_i_1_n_0,counter_reg[2]}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    counter0_carry__0
       (.CI(counter0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_counter0_carry__0_CO_UNCONNECTED[7:5],counter0_carry__0_n_3,counter0_carry__0_n_4,counter0_carry__0_n_5,counter0_carry__0_n_6,counter0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_counter0_carry__0_O_UNCONNECTED[7:6],p_0_in__1[15:10]}),
        .S({1'b0,1'b0,counter_reg[15:10]}));
  LUT1 #(
    .INIT(2'h1)) 
    counter0_carry_i_1
       (.I0(counter_reg[3]),
        .O(counter0_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    \counter[15]_i_1__1 
       (.I0(FRAME_START),
        .I1(frame_start_del),
        .O(START0));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[10] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[10]),
        .Q(counter_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[11] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[11]),
        .Q(counter_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[12] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[12]),
        .Q(counter_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[13] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[13]),
        .Q(counter_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[14] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[14]),
        .Q(counter_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[15] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[15]),
        .Q(counter_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[2] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[2]),
        .Q(counter_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[3] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[3]),
        .Q(counter_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[4] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[4]),
        .Q(counter_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[5] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[5]),
        .Q(counter_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[6] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[6]),
        .Q(counter_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[7] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[7]),
        .Q(counter_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[8] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[8]),
        .Q(counter_reg[8]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[9] 
       (.C(clk_i),
        .CE(START0),
        .CLR(AR),
        .D(p_0_in__1[9]),
        .Q(counter_reg[9]));
  LUT5 #(
    .INIT(32'h2F20202F)) 
    \final_byte_count[10]_i_1 
       (.I0(\final_byte_count_reg[15] [8]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [10]),
        .I4(\final_byte_count_reg[10] ),
        .O(D[8]));
  LUT5 #(
    .INIT(32'h2F20202F)) 
    \final_byte_count[11]_i_1 
       (.I0(\final_byte_count_reg[15] [9]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [11]),
        .I4(\final_byte_count_reg[11] ),
        .O(D[9]));
  LUT6 #(
    .INIT(64'h2F20202F2F202F20)) 
    \final_byte_count[12]_i_1 
       (.I0(\final_byte_count_reg[15] [10]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [12]),
        .I4(\final_byte_count_reg[11] ),
        .I5(\final_byte_count_reg[15]_0 [11]),
        .O(D[10]));
  LUT6 #(
    .INIT(64'h202F2F202F202F20)) 
    \final_byte_count[13]_i_1 
       (.I0(\final_byte_count_reg[15] [11]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [13]),
        .I4(\final_byte_count_reg[13] ),
        .I5(\final_byte_count_reg[15]_0 [12]),
        .O(D[11]));
  LUT5 #(
    .INIT(32'h202F2F20)) 
    \final_byte_count[14]_i_1 
       (.I0(\final_byte_count_reg[15] [12]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [14]),
        .I4(\final_byte_count_reg[14] ),
        .O(D[12]));
  LUT6 #(
    .INIT(64'h202F2F202F202F20)) 
    \final_byte_count[15]_i_1 
       (.I0(\final_byte_count_reg[15] [13]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [15]),
        .I4(\final_byte_count_reg[14] ),
        .I5(\final_byte_count_reg[15]_0 [14]),
        .O(D[13]));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \final_byte_count[15]_i_2 
       (.I0(\final_byte_count[15]_i_4_n_0 ),
        .I1(Q[11]),
        .I2(Q[10]),
        .I3(Q[4]),
        .I4(Q[12]),
        .I5(\final_byte_count[15]_i_5_n_0 ),
        .O(\final_byte_count[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \final_byte_count[15]_i_4 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[5]),
        .I3(Q[13]),
        .I4(Q[2]),
        .I5(Q[3]),
        .O(\final_byte_count[15]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \final_byte_count[15]_i_5 
       (.I0(Q[8]),
        .I1(Q[7]),
        .I2(Q[9]),
        .I3(Q[6]),
        .O(\final_byte_count[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hE0EFEFE0EFE0EFE0)) 
    \final_byte_count[2]_i_1 
       (.I0(\final_byte_count_reg[15] [0]),
        .I1(\final_byte_count[5]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [2]),
        .I4(\final_byte_count_reg[15]_0 [0]),
        .I5(\final_byte_count_reg[15]_0 [1]),
        .O(D[0]));
  LUT5 #(
    .INIT(32'hEFE0E0EF)) 
    \final_byte_count[3]_i_1 
       (.I0(\final_byte_count_reg[15] [1]),
        .I1(\final_byte_count[5]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [3]),
        .I4(\final_byte_count_reg[3] ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'hEFE0E0EF)) 
    \final_byte_count[4]_i_1 
       (.I0(\final_byte_count_reg[15] [2]),
        .I1(\final_byte_count[5]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [4]),
        .I4(\final_byte_count_reg[4] ),
        .O(D[2]));
  LUT5 #(
    .INIT(32'hEFE0E0EF)) 
    \final_byte_count[5]_i_1 
       (.I0(\final_byte_count_reg[15] [3]),
        .I1(\final_byte_count[5]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [5]),
        .I4(\final_byte_count_reg[5] ),
        .O(D[3]));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \final_byte_count[5]_i_2 
       (.I0(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I1(Q[4]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[5]),
        .I5(\final_byte_count[5]_i_4_n_0 ),
        .O(\final_byte_count[5]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair418" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \final_byte_count[5]_i_4 
       (.I0(Q[2]),
        .I1(Q[3]),
        .O(\final_byte_count[5]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h2F20202F)) 
    \final_byte_count[6]_i_1 
       (.I0(\final_byte_count_reg[15] [4]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [6]),
        .I4(\final_byte_count_reg[6] ),
        .O(D[4]));
  LUT6 #(
    .INIT(64'h2F20202F2F202F20)) 
    \final_byte_count[7]_i_1 
       (.I0(\final_byte_count_reg[15] [5]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [7]),
        .I4(\final_byte_count_reg[6] ),
        .I5(\final_byte_count_reg[15]_0 [6]),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h2F20202F)) 
    \final_byte_count[8]_i_1 
       (.I0(\final_byte_count_reg[15] [6]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [8]),
        .I4(\final_byte_count_reg[8] ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h2F20202F)) 
    \final_byte_count[9]_i_1 
       (.I0(\final_byte_count_reg[15] [7]),
        .I1(\final_byte_count[15]_i_2_n_0 ),
        .I2(load_CRC8),
        .I3(\final_byte_count_reg[15]_0 [9]),
        .I4(\final_byte_count_reg[9] ),
        .O(D[7]));
  (* SOFT_HLUTNM = "soft_lutpair410" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[0]_i_1 
       (.I0(\length_register_reg[15] [0]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [16]),
        .O(\TX_DATA_REG_reg[15] [0]));
  (* SOFT_HLUTNM = "soft_lutpair413" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[10]_i_1 
       (.I0(\length_register_reg[15] [10]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [26]),
        .O(\TX_DATA_REG_reg[15] [10]));
  (* SOFT_HLUTNM = "soft_lutpair412" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[11]_i_1 
       (.I0(\length_register_reg[15] [11]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [27]),
        .O(\TX_DATA_REG_reg[15] [11]));
  (* SOFT_HLUTNM = "soft_lutpair411" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[12]_i_1 
       (.I0(\length_register_reg[15] [12]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [28]),
        .O(\TX_DATA_REG_reg[15] [12]));
  (* SOFT_HLUTNM = "soft_lutpair410" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[13]_i_1 
       (.I0(\length_register_reg[15] [13]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [29]),
        .O(\TX_DATA_REG_reg[15] [13]));
  (* SOFT_HLUTNM = "soft_lutpair415" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[14]_i_1 
       (.I0(\length_register_reg[15] [14]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [30]),
        .O(\TX_DATA_REG_reg[15] [14]));
  LUT6 #(
    .INIT(64'h0003002000000000)) 
    \length_register[15]_i_1 
       (.I0(vlan_enabled_int),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(Q[1]),
        .I5(\length_register[15]_i_3_n_0 ),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair417" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[15]_i_2 
       (.I0(\length_register_reg[15] [15]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [31]),
        .O(\TX_DATA_REG_reg[15] [15]));
  (* SOFT_HLUTNM = "soft_lutpair408" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \length_register[15]_i_3 
       (.I0(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I1(Q[5]),
        .I2(Q[4]),
        .O(\length_register[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \length_register[15]_i_4 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(\TX_DATA_VALID_REG[7]_i_3_n_0 ),
        .I3(Q[5]),
        .I4(Q[4]),
        .I5(\length_register[15]_i_5_n_0 ),
        .O(\length_register[15]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair418" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \length_register[15]_i_5 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(vlan_enabled_int),
        .O(\length_register[15]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair411" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[1]_i_1 
       (.I0(\length_register_reg[15] [1]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [17]),
        .O(\TX_DATA_REG_reg[15] [1]));
  (* SOFT_HLUTNM = "soft_lutpair412" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[2]_i_1 
       (.I0(\length_register_reg[15] [2]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [18]),
        .O(\TX_DATA_REG_reg[15] [2]));
  (* SOFT_HLUTNM = "soft_lutpair413" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[3]_i_1 
       (.I0(\length_register_reg[15] [3]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [19]),
        .O(\TX_DATA_REG_reg[15] [3]));
  (* SOFT_HLUTNM = "soft_lutpair414" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[4]_i_1 
       (.I0(\length_register_reg[15] [4]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [20]),
        .O(\TX_DATA_REG_reg[15] [4]));
  (* SOFT_HLUTNM = "soft_lutpair415" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[5]_i_1 
       (.I0(\length_register_reg[15] [5]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [21]),
        .O(\TX_DATA_REG_reg[15] [5]));
  (* SOFT_HLUTNM = "soft_lutpair416" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[6]_i_1 
       (.I0(\length_register_reg[15] [6]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [22]),
        .O(\TX_DATA_REG_reg[15] [6]));
  (* SOFT_HLUTNM = "soft_lutpair417" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[7]_i_1 
       (.I0(\length_register_reg[15] [7]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [23]),
        .O(\TX_DATA_REG_reg[15] [7]));
  (* SOFT_HLUTNM = "soft_lutpair416" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[8]_i_1 
       (.I0(\length_register_reg[15] [8]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [24]),
        .O(\TX_DATA_REG_reg[15] [8]));
  (* SOFT_HLUTNM = "soft_lutpair414" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \length_register[9]_i_1 
       (.I0(\length_register_reg[15] [9]),
        .I1(\length_register[15]_i_4_n_0 ),
        .I2(\length_register_reg[15] [25]),
        .O(\TX_DATA_REG_reg[15] [9]));
endmodule

(* ORIG_REF_NAME = "cfg_crc" *) 
module switch_elements_cfg_crc
   (Q,
    rst_i,
    out,
    \dat_o_reg[0]_0 ,
    clk_i);
  output [4:0]Q;
  input rst_i;
  input out;
  input \dat_o_reg[0]_0 ;
  input clk_i;

  wire [4:0]Q;
  wire clk_i;
  wire \dat_o[0]_i_1__0_n_0 ;
  wire \dat_o[1]_i_1__0_n_0 ;
  wire \dat_o[2]_i_1__0_n_0 ;
  wire \dat_o[3]_i_1__0_n_0 ;
  wire \dat_o[4]_i_1__0_n_0 ;
  wire \dat_o[4]_i_2_n_0 ;
  wire \dat_o_reg[0]_0 ;
  wire out;
  wire rst_i;

  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \dat_o[0]_i_1__0 
       (.I0(\dat_o_reg[0]_0 ),
        .I1(Q[4]),
        .I2(rst_i),
        .O(\dat_o[0]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dat_o[1]_i_1__0 
       (.I0(Q[0]),
        .I1(rst_i),
        .O(\dat_o[1]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \dat_o[2]_i_1__0 
       (.I0(Q[1]),
        .I1(Q[4]),
        .I2(\dat_o_reg[0]_0 ),
        .I3(rst_i),
        .O(\dat_o[2]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dat_o[3]_i_1__0 
       (.I0(Q[2]),
        .I1(rst_i),
        .O(\dat_o[3]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \dat_o[4]_i_1__0 
       (.I0(rst_i),
        .I1(out),
        .O(\dat_o[4]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dat_o[4]_i_2 
       (.I0(Q[3]),
        .I1(rst_i),
        .O(\dat_o[4]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \dat_o_reg[0] 
       (.C(clk_i),
        .CE(\dat_o[4]_i_1__0_n_0 ),
        .CLR(rst_i),
        .D(\dat_o[0]_i_1__0_n_0 ),
        .Q(Q[0]));
  FDCE #(
    .INIT(1'b0)) 
    \dat_o_reg[1] 
       (.C(clk_i),
        .CE(\dat_o[4]_i_1__0_n_0 ),
        .CLR(rst_i),
        .D(\dat_o[1]_i_1__0_n_0 ),
        .Q(Q[1]));
  FDCE #(
    .INIT(1'b0)) 
    \dat_o_reg[2] 
       (.C(clk_i),
        .CE(\dat_o[4]_i_1__0_n_0 ),
        .CLR(rst_i),
        .D(\dat_o[2]_i_1__0_n_0 ),
        .Q(Q[2]));
  FDCE #(
    .INIT(1'b0)) 
    \dat_o_reg[3] 
       (.C(clk_i),
        .CE(\dat_o[4]_i_1__0_n_0 ),
        .CLR(rst_i),
        .D(\dat_o[3]_i_1__0_n_0 ),
        .Q(Q[3]));
  FDCE #(
    .INIT(1'b0)) 
    \dat_o_reg[4] 
       (.C(clk_i),
        .CE(\dat_o[4]_i_1__0_n_0 ),
        .CLR(rst_i),
        .D(\dat_o[4]_i_2_n_0 ),
        .Q(Q[4]));
endmodule

(* ORIG_REF_NAME = "counter" *) 
module switch_elements_counter
   (\value_reg[0]_0 ,
    \value_reg[1]_0 ,
    \value_reg[9]_0 ,
    \value_reg[10]_0 ,
    \value_reg[11]_0 ,
    \value_reg[7]_0 ,
    \value_reg[6]_0 ,
    \value_reg[2]_0 ,
    jumbo_frame0,
    \value_reg[8]_0 ,
    \value_reg[5]_0 ,
    \value_reg[4]_0 ,
    \value_reg[4]_1 ,
    \value_reg[1]_1 ,
    \value_reg[1]_2 ,
    length_256_5110,
    length_512_10230,
    length_65_1270,
    padded_frame0,
    small_error0,
    length_128_2550,
    \value_reg[6]_1 ,
    Q,
    large_error_reg,
    large_error_reg_0,
    get_terminator,
    jumbo_enable,
    large_error_i_4_0,
    \value_reg[9]_1 ,
    tagged_frame,
    vlan_enable,
    clk_i,
    reset_dcm,
    \value_reg[10]_1 ,
    \value_reg[7]_1 ,
    \value_reg[6]_2 ,
    \value_reg[5]_1 ,
    \value_reg[1]_3 ,
    \value_reg[0]_1 );
  output \value_reg[0]_0 ;
  output \value_reg[1]_0 ;
  output \value_reg[9]_0 ;
  output \value_reg[10]_0 ;
  output \value_reg[11]_0 ;
  output \value_reg[7]_0 ;
  output \value_reg[6]_0 ;
  output \value_reg[2]_0 ;
  output jumbo_frame0;
  output \value_reg[8]_0 ;
  output \value_reg[5]_0 ;
  output \value_reg[4]_0 ;
  output \value_reg[4]_1 ;
  output \value_reg[1]_1 ;
  output \value_reg[1]_2 ;
  output length_256_5110;
  output length_512_10230;
  output length_65_1270;
  output padded_frame0;
  output small_error0;
  output length_128_2550;
  output \value_reg[6]_1 ;
  input [2:0]Q;
  input large_error_reg;
  input large_error_reg_0;
  input get_terminator;
  input jumbo_enable;
  input [0:0]large_error_i_4_0;
  input \value_reg[9]_1 ;
  input tagged_frame;
  input vlan_enable;
  input clk_i;
  input reset_dcm;
  input \value_reg[10]_1 ;
  input \value_reg[7]_1 ;
  input \value_reg[6]_2 ;
  input \value_reg[5]_1 ;
  input [0:0]\value_reg[1]_3 ;
  input \value_reg[0]_1 ;

  wire [2:0]Q;
  wire clk_i;
  wire [11:2]frame_cnt;
  wire get_terminator;
  wire jumbo_enable;
  wire jumbo_frame0;
  wire jumbo_frame_i_2_n_0;
  wire jumbo_frame_i_3_n_0;
  wire jumbo_frame_i_4_n_0;
  wire large_error_i_3_n_0;
  wire [0:0]large_error_i_4_0;
  wire large_error_i_4_n_0;
  wire large_error_i_5_n_0;
  wire large_error_i_7_n_0;
  wire large_error_i_9_n_0;
  wire large_error_reg;
  wire large_error_reg_0;
  wire length_128_2550;
  wire length_128_255_i_2_n_0;
  wire length_256_5110;
  wire length_256_511_i_2_n_0;
  wire length_512_10230;
  wire length_65_1270;
  wire length_65_127_i_2_n_0;
  wire length_65_127_i_3_n_0;
  wire [11:2]p_0_in;
  wire padded_frame0;
  wire padded_frame_i_2_n_0;
  wire reset_dcm;
  wire small_error0;
  wire small_error_i_2_n_0;
  wire tagged_frame;
  wire \value[3]_i_1_n_0 ;
  wire \value[4]_i_1_n_0 ;
  wire \value[8]_i_1_n_0 ;
  wire \value[9]_i_1_n_0 ;
  wire \value_reg[0]_0 ;
  wire \value_reg[0]_1 ;
  wire \value_reg[10]_0 ;
  wire \value_reg[10]_1 ;
  wire \value_reg[11]_0 ;
  wire \value_reg[1]_0 ;
  wire \value_reg[1]_1 ;
  wire \value_reg[1]_2 ;
  wire [0:0]\value_reg[1]_3 ;
  wire \value_reg[2]_0 ;
  wire \value_reg[4]_0 ;
  wire \value_reg[4]_1 ;
  wire \value_reg[5]_0 ;
  wire \value_reg[5]_1 ;
  wire \value_reg[6]_0 ;
  wire \value_reg[6]_1 ;
  wire \value_reg[6]_2 ;
  wire \value_reg[7]_0 ;
  wire \value_reg[7]_1 ;
  wire \value_reg[8]_0 ;
  wire \value_reg[9]_0 ;
  wire \value_reg[9]_1 ;
  wire vlan_enable;

  LUT6 #(
    .INIT(64'h0080008000808080)) 
    jumbo_frame_i_1
       (.I0(large_error_i_3_n_0),
        .I1(get_terminator),
        .I2(jumbo_enable),
        .I3(jumbo_frame_i_2_n_0),
        .I4(jumbo_frame_i_3_n_0),
        .I5(jumbo_frame_i_4_n_0),
        .O(jumbo_frame0));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'hE)) 
    jumbo_frame_i_2
       (.I0(\value_reg[10]_0 ),
        .I1(frame_cnt[11]),
        .O(jumbo_frame_i_2_n_0));
  LUT6 #(
    .INIT(64'h8888888088808880)) 
    jumbo_frame_i_3
       (.I0(\value_reg[6]_0 ),
        .I1(\value_reg[5]_0 ),
        .I2(frame_cnt[3]),
        .I3(\value_reg[4]_0 ),
        .I4(\value_reg[1]_0 ),
        .I5(frame_cnt[2]),
        .O(jumbo_frame_i_3_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    jumbo_frame_i_4
       (.I0(frame_cnt[8]),
        .I1(\value_reg[7]_0 ),
        .I2(frame_cnt[11]),
        .I3(frame_cnt[9]),
        .O(jumbo_frame_i_4_n_0));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFFFFFF4)) 
    large_error_i_1
       (.I0(large_error_reg),
        .I1(large_error_i_3_n_0),
        .I2(large_error_i_4_n_0),
        .I3(frame_cnt[11]),
        .I4(\value_reg[10]_0 ),
        .I5(large_error_i_5_n_0),
        .O(\value_reg[11]_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    large_error_i_10
       (.I0(\value_reg[4]_0 ),
        .I1(\value_reg[5]_0 ),
        .O(\value_reg[4]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h7)) 
    large_error_i_11
       (.I0(\value_reg[1]_0 ),
        .I1(frame_cnt[2]),
        .O(\value_reg[1]_2 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    large_error_i_3
       (.I0(\value_reg[2]_0 ),
        .I1(\value_reg[6]_0 ),
        .I2(\value_reg[7]_0 ),
        .I3(\value_reg[8]_0 ),
        .O(large_error_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    large_error_i_4
       (.I0(large_error_i_7_n_0),
        .I1(large_error_reg_0),
        .I2(\value_reg[7]_0 ),
        .I3(\value_reg[6]_0 ),
        .I4(frame_cnt[3]),
        .I5(\value_reg[0]_0 ),
        .O(large_error_i_4_n_0));
  LUT6 #(
    .INIT(64'h00000000777F7777)) 
    large_error_i_5
       (.I0(\value_reg[5]_0 ),
        .I1(\value_reg[6]_0 ),
        .I2(\value_reg[4]_0 ),
        .I3(frame_cnt[3]),
        .I4(large_error_i_9_n_0),
        .I5(jumbo_frame_i_4_n_0),
        .O(large_error_i_5_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    large_error_i_6
       (.I0(\value_reg[6]_0 ),
        .I1(tagged_frame),
        .I2(vlan_enable),
        .O(\value_reg[6]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    large_error_i_7
       (.I0(large_error_i_4_0),
        .I1(frame_cnt[9]),
        .I2(frame_cnt[11]),
        .I3(\value_reg[10]_0 ),
        .I4(frame_cnt[8]),
        .O(large_error_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    large_error_i_9
       (.I0(frame_cnt[2]),
        .I1(\value_reg[1]_0 ),
        .I2(\value_reg[0]_0 ),
        .O(large_error_i_9_n_0));
  LUT5 #(
    .INIT(32'h0000E000)) 
    length_128_255_i_1
       (.I0(\value_reg[6]_0 ),
        .I1(length_128_255_i_2_n_0),
        .I2(\value_reg[7]_0 ),
        .I3(get_terminator),
        .I4(\value_reg[8]_0 ),
        .O(length_128_2550));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    length_128_255_i_2
       (.I0(\value_reg[0]_0 ),
        .I1(\value_reg[1]_0 ),
        .I2(frame_cnt[2]),
        .I3(frame_cnt[3]),
        .I4(\value_reg[4]_0 ),
        .I5(\value_reg[5]_0 ),
        .O(length_128_255_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    length_128_255_i_3
       (.I0(frame_cnt[8]),
        .I1(\value_reg[10]_0 ),
        .I2(frame_cnt[11]),
        .I3(frame_cnt[9]),
        .O(\value_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    length_256_511_i_1
       (.I0(length_256_511_i_2_n_0),
        .I1(frame_cnt[8]),
        .I2(frame_cnt[9]),
        .I3(get_terminator),
        .I4(\value_reg[10]_0 ),
        .I5(frame_cnt[11]),
        .O(length_256_5110));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    length_256_511_i_2
       (.I0(\value_reg[7]_0 ),
        .I1(\value_reg[6]_0 ),
        .I2(\value_reg[5]_0 ),
        .I3(\value_reg[4]_0 ),
        .I4(frame_cnt[3]),
        .I5(length_65_127_i_3_n_0),
        .O(length_256_511_i_2_n_0));
  LUT6 #(
    .INIT(64'h000000E000000000)) 
    length_512_1023_i_1
       (.I0(length_256_511_i_2_n_0),
        .I1(frame_cnt[8]),
        .I2(frame_cnt[9]),
        .I3(frame_cnt[11]),
        .I4(\value_reg[10]_0 ),
        .I5(get_terminator),
        .O(length_512_10230));
  LUT6 #(
    .INIT(64'h1011101011111111)) 
    length_65_127_i_1
       (.I0(length_65_127_i_2_n_0),
        .I1(\value_reg[7]_0 ),
        .I2(\value_reg[6]_0 ),
        .I3(length_65_127_i_3_n_0),
        .I4(frame_cnt[3]),
        .I5(small_error_i_2_n_0),
        .O(length_65_1270));
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    length_65_127_i_2
       (.I0(frame_cnt[9]),
        .I1(frame_cnt[11]),
        .I2(\value_reg[10]_0 ),
        .I3(frame_cnt[8]),
        .I4(get_terminator),
        .O(length_65_127_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'h01)) 
    length_65_127_i_3
       (.I0(frame_cnt[2]),
        .I1(\value_reg[1]_0 ),
        .I2(\value_reg[0]_0 ),
        .O(length_65_127_i_3_n_0));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT5 #(
    .INIT(32'h00020000)) 
    padded_frame_i_1
       (.I0(padded_frame_i_2_n_0),
        .I1(frame_cnt[2]),
        .I2(\value_reg[1]_0 ),
        .I3(\value_reg[0]_0 ),
        .I4(frame_cnt[3]),
        .O(padded_frame0));
  LUT5 #(
    .INIT(32'h00000020)) 
    padded_frame_i_2
       (.I0(small_error_i_2_n_0),
        .I1(frame_cnt[8]),
        .I2(get_terminator),
        .I3(\value_reg[6]_0 ),
        .I4(\value_reg[7]_0 ),
        .O(padded_frame_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    small_error_i_1
       (.I0(\value_reg[7]_0 ),
        .I1(\value_reg[6]_0 ),
        .I2(get_terminator),
        .I3(frame_cnt[8]),
        .I4(small_error_i_2_n_0),
        .I5(frame_cnt[3]),
        .O(small_error0));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    small_error_i_2
       (.I0(\value_reg[10]_0 ),
        .I1(frame_cnt[11]),
        .I2(frame_cnt[9]),
        .I3(\value_reg[5]_0 ),
        .I4(\value_reg[4]_0 ),
        .O(small_error_i_2_n_0));
  LUT6 #(
    .INIT(64'h7878787878787800)) 
    \value[11]_i_1 
       (.I0(\value_reg[9]_0 ),
        .I1(\value_reg[10]_0 ),
        .I2(frame_cnt[11]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(p_0_in[11]));
  LUT5 #(
    .INIT(32'h00800000)) 
    \value[11]_i_2 
       (.I0(frame_cnt[9]),
        .I1(frame_cnt[8]),
        .I2(\value_reg[6]_0 ),
        .I3(\value_reg[2]_0 ),
        .I4(\value_reg[7]_0 ),
        .O(\value_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h7878787878787800)) 
    \value[2]_i_1 
       (.I0(\value_reg[0]_0 ),
        .I1(\value_reg[1]_0 ),
        .I2(frame_cnt[2]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(p_0_in[2]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT5 #(
    .INIT(32'h15554000)) 
    \value[3]_i_1 
       (.I0(\value_reg[9]_1 ),
        .I1(frame_cnt[2]),
        .I2(\value_reg[1]_0 ),
        .I3(\value_reg[0]_0 ),
        .I4(frame_cnt[3]),
        .O(\value[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    \value[4]_i_1 
       (.I0(\value_reg[9]_1 ),
        .I1(\value_reg[1]_0 ),
        .I2(\value_reg[0]_0 ),
        .I3(frame_cnt[3]),
        .I4(frame_cnt[2]),
        .I5(\value_reg[4]_0 ),
        .O(\value[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \value[5]_i_2 
       (.I0(\value_reg[1]_0 ),
        .I1(\value_reg[0]_0 ),
        .I2(frame_cnt[3]),
        .I3(frame_cnt[2]),
        .O(\value_reg[1]_1 ));
  LUT5 #(
    .INIT(32'h51550400)) 
    \value[8]_i_1 
       (.I0(\value_reg[9]_1 ),
        .I1(\value_reg[6]_0 ),
        .I2(\value_reg[2]_0 ),
        .I3(\value_reg[7]_0 ),
        .I4(frame_cnt[8]),
        .O(\value[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5155555504000000)) 
    \value[9]_i_1 
       (.I0(\value_reg[9]_1 ),
        .I1(\value_reg[7]_0 ),
        .I2(\value_reg[2]_0 ),
        .I3(\value_reg[6]_0 ),
        .I4(frame_cnt[8]),
        .I5(frame_cnt[9]),
        .O(\value[9]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \value[9]_i_2 
       (.I0(frame_cnt[2]),
        .I1(frame_cnt[3]),
        .I2(\value_reg[0]_0 ),
        .I3(\value_reg[1]_0 ),
        .I4(\value_reg[5]_0 ),
        .I5(\value_reg[4]_0 ),
        .O(\value_reg[2]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value_reg[0]_1 ),
        .Q(\value_reg[0]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value_reg[10]_1 ),
        .Q(\value_reg[10]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_0_in[11]),
        .Q(frame_cnt[11]));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value_reg[1]_3 ),
        .Q(\value_reg[1]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(p_0_in[2]),
        .Q(frame_cnt[2]));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value[3]_i_1_n_0 ),
        .Q(frame_cnt[3]));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value[4]_i_1_n_0 ),
        .Q(\value_reg[4]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value_reg[5]_1 ),
        .Q(\value_reg[5]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value_reg[6]_2 ),
        .Q(\value_reg[6]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value_reg[7]_1 ),
        .Q(\value_reg[7]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value[8]_i_1_n_0 ),
        .Q(frame_cnt[8]));
  FDCE #(
    .INIT(1'b0)) 
    \value_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\value[9]_i_1_n_0 ),
        .Q(frame_cnt[9]));
endmodule

(* ORIG_REF_NAME = "decode" *) 
module switch_elements_decode
   (ready_o,
    Q,
    \index_reg[4]_0 ,
    \FSM_sequential_state_reg[0]_0 ,
    \FSM_sequential_state_reg[2]_0 ,
    \FSM_sequential_state_reg[1]_0 ,
    q_o,
    clk_i,
    rst_i,
    md16_nd,
    \FSM_sequential_state_reg[2]_1 ,
    \FSM_sequential_state_reg[2]_2 ,
    \FSM_sequential_state_reg[0]_1 ,
    CO,
    \FSM_sequential_state_reg[0]_2 ,
    \FSM_sequential_state_reg[0]_3 ,
    D);
  output ready_o;
  output [0:0]Q;
  output \index_reg[4]_0 ;
  output \FSM_sequential_state_reg[0]_0 ;
  output \FSM_sequential_state_reg[2]_0 ;
  output \FSM_sequential_state_reg[1]_0 ;
  output [3:0]q_o;
  input clk_i;
  input rst_i;
  input md16_nd;
  input \FSM_sequential_state_reg[2]_1 ;
  input \FSM_sequential_state_reg[2]_2 ;
  input \FSM_sequential_state_reg[0]_1 ;
  input [0:0]CO;
  input [0:0]\FSM_sequential_state_reg[0]_2 ;
  input [0:0]\FSM_sequential_state_reg[0]_3 ;
  input [0:0]D;

  wire [0:0]CO;
  wire [0:0]D;
  wire \FSM_sequential_state[0]_i_1__0_n_0 ;
  wire \FSM_sequential_state[0]_i_2_n_0 ;
  wire \FSM_sequential_state[2]_i_1_n_0 ;
  wire \FSM_sequential_state[2]_i_3_n_0 ;
  wire \FSM_sequential_state_reg[0]_0 ;
  wire \FSM_sequential_state_reg[0]_1 ;
  wire [0:0]\FSM_sequential_state_reg[0]_2 ;
  wire [0:0]\FSM_sequential_state_reg[0]_3 ;
  wire \FSM_sequential_state_reg[1]_0 ;
  wire \FSM_sequential_state_reg[2]_0 ;
  wire \FSM_sequential_state_reg[2]_1 ;
  wire \FSM_sequential_state_reg[2]_2 ;
  wire [0:0]Q;
  wire clk_i;
  wire [4:0]index;
  wire \index[0]_i_1_n_0 ;
  wire \index[1]_i_1_n_0 ;
  wire \index[1]_i_2_n_0 ;
  wire \index[2]_i_1_n_0 ;
  wire \index[2]_i_2_n_0 ;
  wire \index[3]_i_1_n_0 ;
  wire \index[3]_i_2_n_0 ;
  wire \index[4]_i_2_n_0 ;
  wire \index[4]_i_3_n_0 ;
  wire \index[4]_i_4_n_0 ;
  wire \index_reg[4]_0 ;
  wire md16_nd;
  wire nd_o_buff;
  wire nd_o_buff_i_1_n_0;
  wire [1:0]p_0_in;
  wire [1:0]p_1_in;
  wire [3:0]p_3_out;
  wire [3:0]q_o;
  wire ready_o;
  wire rst_i;
  wire [2:1]state;
  wire \str_buffer[0]_i_1_n_0 ;
  wire \str_buffer[0]_i_2_n_0 ;
  wire \str_buffer[0]_i_3_n_0 ;
  wire \str_buffer[0]_i_4_n_0 ;
  wire \str_buffer[1]_i_1_n_0 ;
  wire \str_buffer[1]_i_2_n_0 ;
  wire \str_buffer[1]_i_3_n_0 ;
  wire \str_buffer[1]_i_4_n_0 ;
  wire \str_buffer[1]_i_5_n_0 ;
  wire \str_buffer[1]_i_6_n_0 ;
  wire \str_buffer[2]_i_1_n_0 ;
  wire \str_buffer[2]_i_2_n_0 ;
  wire \str_buffer[3]_i_1_n_0 ;
  wire \str_buffer[3]_i_2_n_0 ;
  wire \str_buffer[3]_i_3_n_0 ;
  wire \str_buffer[4]_i_1_n_0 ;
  wire \str_buffer[4]_i_2_n_0 ;
  wire \str_buffer[4]_i_3_n_0 ;
  wire \str_buffer[5]_i_1_n_0 ;
  wire \str_buffer[5]_i_2_n_0 ;
  wire \str_buffer[5]_i_3_n_0 ;
  wire \str_buffer[5]_i_4_n_0 ;
  wire \str_buffer[6]_i_1_n_0 ;
  wire \str_buffer[6]_i_2_n_0 ;
  wire \str_buffer[6]_i_3_n_0 ;
  wire \str_buffer[6]_i_4_n_0 ;
  wire \str_buffer[7]_i_1_n_0 ;
  wire \str_buffer[7]_i_2_n_0 ;
  wire \str_buffer[7]_i_3_n_0 ;
  wire \str_buffer[7]_i_4_n_0 ;
  wire \str_buffer[7]_i_5_n_0 ;
  wire \str_buffer_reg_n_0_[0] ;
  wire \str_buffer_reg_n_0_[1] ;
  wire \str_buffer_reg_n_0_[2] ;
  wire \str_buffer_reg_n_0_[3] ;

  LUT6 #(
    .INIT(64'h80808080808080F0)) 
    \FSM_sequential_state[0]_i_1__0 
       (.I0(\FSM_sequential_state[0]_i_2_n_0 ),
        .I1(\FSM_sequential_state_reg[0]_1 ),
        .I2(\index_reg[4]_0 ),
        .I3(state[2]),
        .I4(state[1]),
        .I5(Q),
        .O(\FSM_sequential_state[0]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h001D1D1D35000000)) 
    \FSM_sequential_state[0]_i_2 
       (.I0(Q),
        .I1(state[1]),
        .I2(state[2]),
        .I3(CO),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\FSM_sequential_state_reg[0]_3 ),
        .O(\FSM_sequential_state[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_state[1]_i_5__0 
       (.I0(state[1]),
        .I1(state[2]),
        .O(\FSM_sequential_state_reg[1]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'h74)) 
    \FSM_sequential_state[1]_i_6__0 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(Q),
        .O(\FSM_sequential_state_reg[2]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'h34)) 
    \FSM_sequential_state[1]_i_7__0 
       (.I0(Q),
        .I1(state[2]),
        .I2(state[1]),
        .O(\FSM_sequential_state_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0A8008A000800880)) 
    \FSM_sequential_state[2]_i_1 
       (.I0(\FSM_sequential_state[2]_i_3_n_0 ),
        .I1(\FSM_sequential_state_reg[2]_1 ),
        .I2(state[2]),
        .I3(state[1]),
        .I4(Q),
        .I5(\FSM_sequential_state_reg[2]_2 ),
        .O(\FSM_sequential_state[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \FSM_sequential_state[2]_i_3 
       (.I0(index[0]),
        .I1(index[3]),
        .I2(index[2]),
        .I3(index[1]),
        .I4(index[4]),
        .I5(\FSM_sequential_state_reg[0]_3 ),
        .O(\FSM_sequential_state[2]_i_3_n_0 ));
  (* FSM_ENCODED_STATES = "pause:001,one_1:010,reset:000,two_0:011,one_0:101,two_1:100" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[0] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\FSM_sequential_state[0]_i_1__0_n_0 ),
        .Q(Q));
  (* FSM_ENCODED_STATES = "pause:001,one_1:010,reset:000,two_0:011,one_0:101,two_1:100" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[1] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(D),
        .Q(state[1]));
  (* FSM_ENCODED_STATES = "pause:001,one_1:010,reset:000,two_0:011,one_0:101,two_1:100" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[2] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\FSM_sequential_state[2]_i_1_n_0 ),
        .Q(state[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \decoded_o[0]_i_1 
       (.I0(p_0_in[0]),
        .I1(p_0_in[1]),
        .O(p_3_out[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \decoded_o[1]_i_1 
       (.I0(p_1_in[0]),
        .I1(p_1_in[1]),
        .O(p_3_out[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \decoded_o[2]_i_1 
       (.I0(\str_buffer_reg_n_0_[2] ),
        .I1(\str_buffer_reg_n_0_[3] ),
        .O(p_3_out[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \decoded_o[3]_i_1 
       (.I0(\str_buffer_reg_n_0_[0] ),
        .I1(\str_buffer_reg_n_0_[1] ),
        .O(p_3_out[3]));
  FDCE #(
    .INIT(1'b0)) 
    \decoded_o_reg[0] 
       (.C(clk_i),
        .CE(nd_o_buff),
        .CLR(rst_i),
        .D(p_3_out[0]),
        .Q(q_o[0]));
  FDCE #(
    .INIT(1'b0)) 
    \decoded_o_reg[1] 
       (.C(clk_i),
        .CE(nd_o_buff),
        .CLR(rst_i),
        .D(p_3_out[1]),
        .Q(q_o[1]));
  FDCE #(
    .INIT(1'b0)) 
    \decoded_o_reg[2] 
       (.C(clk_i),
        .CE(nd_o_buff),
        .CLR(rst_i),
        .D(p_3_out[2]),
        .Q(q_o[2]));
  FDCE #(
    .INIT(1'b0)) 
    \decoded_o_reg[3] 
       (.C(clk_i),
        .CE(nd_o_buff),
        .CLR(rst_i),
        .D(p_3_out[3]),
        .Q(q_o[3]));
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT5 #(
    .INIT(32'hF01441F0)) 
    \index[0]_i_1 
       (.I0(index[4]),
        .I1(Q),
        .I2(index[0]),
        .I3(state[1]),
        .I4(state[2]),
        .O(\index[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT4 #(
    .INIT(16'hA0AC)) 
    \index[1]_i_1 
       (.I0(\index[3]_i_2_n_0 ),
        .I1(\index[1]_i_2_n_0 ),
        .I2(index[1]),
        .I3(index[4]),
        .O(\index[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000FE0F0FFE0000)) 
    \index[1]_i_2 
       (.I0(index[3]),
        .I1(index[2]),
        .I2(index[0]),
        .I3(Q),
        .I4(state[2]),
        .I5(state[1]),
        .O(\index[1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT5 #(
    .INIT(32'hFFAAAEAA)) 
    \index[2]_i_1 
       (.I0(\index[2]_i_2_n_0 ),
        .I1(index[1]),
        .I2(index[4]),
        .I3(index[2]),
        .I4(\index[3]_i_2_n_0 ),
        .O(\index[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000C3000000BE0)) 
    \index[2]_i_2 
       (.I0(index[3]),
        .I1(Q),
        .I2(state[2]),
        .I3(state[1]),
        .I4(\str_buffer[1]_i_3_n_0 ),
        .I5(index[0]),
        .O(\index[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAAABBBAAAAA)) 
    \index[3]_i_1 
       (.I0(\index[4]_i_3_n_0 ),
        .I1(index[4]),
        .I2(index[2]),
        .I3(index[1]),
        .I4(index[3]),
        .I5(\index[3]_i_2_n_0 ),
        .O(\index[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT5 #(
    .INIT(32'hFF0408FF)) 
    \index[3]_i_2 
       (.I0(Q),
        .I1(index[0]),
        .I2(index[4]),
        .I3(state[2]),
        .I4(state[1]),
        .O(\index[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \index[4]_i_1 
       (.I0(index[4]),
        .I1(index[1]),
        .I2(index[2]),
        .I3(index[3]),
        .I4(index[0]),
        .O(\index_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFAAAEAEEAEAFFAA)) 
    \index[4]_i_2 
       (.I0(\index[4]_i_3_n_0 ),
        .I1(\index[4]_i_4_n_0 ),
        .I2(Q),
        .I3(index[4]),
        .I4(state[1]),
        .I5(state[2]),
        .O(\index[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000100101100000)) 
    \index[4]_i_3 
       (.I0(\str_buffer[1]_i_3_n_0 ),
        .I1(index[3]),
        .I2(index[0]),
        .I3(Q),
        .I4(state[2]),
        .I5(state[1]),
        .O(\index[4]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT4 #(
    .INIT(16'h4440)) 
    \index[4]_i_4 
       (.I0(index[4]),
        .I1(index[3]),
        .I2(index[2]),
        .I3(index[1]),
        .O(\index[4]_i_4_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \index_reg[0] 
       (.C(md16_nd),
        .CE(\index_reg[4]_0 ),
        .D(\index[0]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(index[0]));
  FDCE #(
    .INIT(1'b0)) 
    \index_reg[1] 
       (.C(md16_nd),
        .CE(\index_reg[4]_0 ),
        .CLR(rst_i),
        .D(\index[1]_i_1_n_0 ),
        .Q(index[1]));
  FDCE #(
    .INIT(1'b0)) 
    \index_reg[2] 
       (.C(md16_nd),
        .CE(\index_reg[4]_0 ),
        .CLR(rst_i),
        .D(\index[2]_i_1_n_0 ),
        .Q(index[2]));
  FDPE #(
    .INIT(1'b1)) 
    \index_reg[3] 
       (.C(md16_nd),
        .CE(\index_reg[4]_0 ),
        .D(\index[3]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(index[3]));
  FDCE #(
    .INIT(1'b0)) 
    \index_reg[4] 
       (.C(md16_nd),
        .CE(\index_reg[4]_0 ),
        .CLR(rst_i),
        .D(\index[4]_i_2_n_0 ),
        .Q(index[4]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAB)) 
    nd_o_buff_i_1
       (.I0(nd_o_buff),
        .I1(index[0]),
        .I2(index[3]),
        .I3(index[2]),
        .I4(index[1]),
        .I5(index[4]),
        .O(nd_o_buff_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    nd_o_buff_reg
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(nd_o_buff_i_1_n_0),
        .Q(nd_o_buff));
  FDCE #(
    .INIT(1'b0)) 
    nd_o_reg
       (.C(clk_i),
        .CE(nd_o_buff),
        .CLR(rst_i),
        .D(nd_o_buff),
        .Q(ready_o));
  LUT5 #(
    .INIT(32'hBBBA888A)) 
    \str_buffer[0]_i_1 
       (.I0(\str_buffer[0]_i_2_n_0 ),
        .I1(\str_buffer[0]_i_3_n_0 ),
        .I2(nd_o_buff),
        .I3(\index_reg[4]_0 ),
        .I4(\str_buffer_reg_n_0_[0] ),
        .O(\str_buffer[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h003C002C002C003C)) 
    \str_buffer[0]_i_2 
       (.I0(index[4]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(Q),
        .I4(index[3]),
        .I5(\str_buffer[0]_i_4_n_0 ),
        .O(\str_buffer[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \str_buffer[0]_i_3 
       (.I0(index[2]),
        .I1(index[1]),
        .I2(index[4]),
        .I3(nd_o_buff),
        .I4(index[3]),
        .I5(\str_buffer[5]_i_4_n_0 ),
        .O(\str_buffer[0]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \str_buffer[0]_i_4 
       (.I0(index[1]),
        .I1(index[2]),
        .O(\str_buffer[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAFFEFAAAA0020)) 
    \str_buffer[1]_i_1 
       (.I0(\str_buffer[1]_i_2_n_0 ),
        .I1(\str_buffer[1]_i_3_n_0 ),
        .I2(\str_buffer[1]_i_4_n_0 ),
        .I3(nd_o_buff),
        .I4(\str_buffer[1]_i_5_n_0 ),
        .I5(\str_buffer_reg_n_0_[1] ),
        .O(\str_buffer[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCCCCCDFCCCC)) 
    \str_buffer[1]_i_2 
       (.I0(index[0]),
        .I1(\str_buffer[7]_i_5_n_0 ),
        .I2(index[1]),
        .I3(index[2]),
        .I4(\str_buffer[6]_i_2_n_0 ),
        .I5(index[3]),
        .O(\str_buffer[1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \str_buffer[1]_i_3 
       (.I0(index[2]),
        .I1(index[1]),
        .I2(index[4]),
        .O(\str_buffer[1]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \str_buffer[1]_i_4 
       (.I0(index[0]),
        .I1(index[3]),
        .O(\str_buffer[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \str_buffer[1]_i_5 
       (.I0(\str_buffer[1]_i_6_n_0 ),
        .I1(index[2]),
        .I2(nd_o_buff),
        .I3(index[4]),
        .I4(index[1]),
        .I5(\str_buffer[5]_i_4_n_0 ),
        .O(\str_buffer[1]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \str_buffer[1]_i_6 
       (.I0(index[0]),
        .I1(index[3]),
        .O(\str_buffer[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFFF00800000)) 
    \str_buffer[2]_i_1 
       (.I0(\str_buffer[2]_i_2_n_0 ),
        .I1(\str_buffer[7]_i_4_n_0 ),
        .I2(index[1]),
        .I3(index[2]),
        .I4(\str_buffer[6]_i_4_n_0 ),
        .I5(\str_buffer_reg_n_0_[2] ),
        .O(\str_buffer[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFCECFCECCCECCCFC)) 
    \str_buffer[2]_i_2 
       (.I0(index[1]),
        .I1(\str_buffer[4]_i_3_n_0 ),
        .I2(\str_buffer[6]_i_2_n_0 ),
        .I3(index[2]),
        .I4(index[0]),
        .I5(index[3]),
        .O(\str_buffer[2]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \str_buffer[3]_i_1 
       (.I0(\str_buffer[3]_i_2_n_0 ),
        .I1(\str_buffer[3]_i_3_n_0 ),
        .I2(\str_buffer_reg_n_0_[3] ),
        .O(\str_buffer[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAFAAAAAAAAABABA)) 
    \str_buffer[3]_i_2 
       (.I0(\str_buffer[7]_i_5_n_0 ),
        .I1(index[3]),
        .I2(\str_buffer[6]_i_2_n_0 ),
        .I3(index[2]),
        .I4(index[1]),
        .I5(index[0]),
        .O(\str_buffer[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000C0000000080)) 
    \str_buffer[3]_i_3 
       (.I0(\str_buffer[5]_i_4_n_0 ),
        .I1(\str_buffer[7]_i_4_n_0 ),
        .I2(index[2]),
        .I3(index[1]),
        .I4(index[3]),
        .I5(index[0]),
        .O(\str_buffer[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFFF00800000)) 
    \str_buffer[4]_i_1 
       (.I0(\str_buffer[4]_i_2_n_0 ),
        .I1(\str_buffer[7]_i_4_n_0 ),
        .I2(index[2]),
        .I3(index[1]),
        .I4(\str_buffer[6]_i_4_n_0 ),
        .I5(p_1_in[0]),
        .O(\str_buffer[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFEFECECFCCCCCCCC)) 
    \str_buffer[4]_i_2 
       (.I0(index[2]),
        .I1(\str_buffer[4]_i_3_n_0 ),
        .I2(index[1]),
        .I3(index[0]),
        .I4(index[3]),
        .I5(\str_buffer[6]_i_2_n_0 ),
        .O(\str_buffer[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT4 #(
    .INIT(16'h002C)) 
    \str_buffer[4]_i_3 
       (.I0(index[4]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(Q),
        .O(\str_buffer[4]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \str_buffer[5]_i_1 
       (.I0(\str_buffer[5]_i_2_n_0 ),
        .I1(\str_buffer[5]_i_3_n_0 ),
        .I2(p_1_in[1]),
        .O(\str_buffer[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCFCCCFCCCCCDC)) 
    \str_buffer[5]_i_2 
       (.I0(index[3]),
        .I1(\str_buffer[7]_i_5_n_0 ),
        .I2(\str_buffer[6]_i_2_n_0 ),
        .I3(index[2]),
        .I4(index[1]),
        .I5(index[0]),
        .O(\str_buffer[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000C0000008000)) 
    \str_buffer[5]_i_3 
       (.I0(\str_buffer[5]_i_4_n_0 ),
        .I1(\str_buffer[7]_i_4_n_0 ),
        .I2(index[1]),
        .I3(index[2]),
        .I4(index[3]),
        .I5(index[0]),
        .O(\str_buffer[5]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'h18)) 
    \str_buffer[5]_i_4 
       (.I0(Q),
        .I1(state[1]),
        .I2(state[2]),
        .O(\str_buffer[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFFFFFE0000000)) 
    \str_buffer[6]_i_1 
       (.I0(\str_buffer[6]_i_2_n_0 ),
        .I1(\str_buffer[6]_i_3_n_0 ),
        .I2(\str_buffer[7]_i_3_n_0 ),
        .I3(\str_buffer[7]_i_4_n_0 ),
        .I4(\str_buffer[6]_i_4_n_0 ),
        .I5(p_0_in[0]),
        .O(\str_buffer[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \str_buffer[6]_i_2 
       (.I0(state[1]),
        .I1(state[2]),
        .I2(Q),
        .O(\str_buffer[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000010)) 
    \str_buffer[6]_i_3 
       (.I0(index[0]),
        .I1(index[3]),
        .I2(\str_buffer[6]_i_2_n_0 ),
        .I3(index[2]),
        .I4(index[1]),
        .I5(\str_buffer[7]_i_5_n_0 ),
        .O(\str_buffer[6]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT5 #(
    .INIT(32'h001800FF)) 
    \str_buffer[6]_i_4 
       (.I0(Q),
        .I1(state[1]),
        .I2(state[2]),
        .I3(index[3]),
        .I4(index[0]),
        .O(\str_buffer[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFFF00800000)) 
    \str_buffer[7]_i_1 
       (.I0(\str_buffer[7]_i_2_n_0 ),
        .I1(\str_buffer[7]_i_3_n_0 ),
        .I2(\str_buffer[7]_i_4_n_0 ),
        .I3(index[3]),
        .I4(index[0]),
        .I5(p_0_in[1]),
        .O(\str_buffer[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT5 #(
    .INIT(32'hEAAAAAAE)) 
    \str_buffer[7]_i_2 
       (.I0(\str_buffer[7]_i_5_n_0 ),
        .I1(\str_buffer[6]_i_2_n_0 ),
        .I2(index[2]),
        .I3(index[1]),
        .I4(index[0]),
        .O(\str_buffer[7]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \str_buffer[7]_i_3 
       (.I0(index[1]),
        .I1(index[2]),
        .O(\str_buffer[7]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \str_buffer[7]_i_4 
       (.I0(index[4]),
        .I1(nd_o_buff),
        .O(\str_buffer[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000F0F00000F0800)) 
    \str_buffer[7]_i_5 
       (.I0(\str_buffer[0]_i_4_n_0 ),
        .I1(index[3]),
        .I2(Q),
        .I3(state[2]),
        .I4(state[1]),
        .I5(index[4]),
        .O(\str_buffer[7]_i_5_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[0] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[0]_i_1_n_0 ),
        .Q(\str_buffer_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[1] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[1]_i_1_n_0 ),
        .Q(\str_buffer_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[2] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[2]_i_1_n_0 ),
        .Q(\str_buffer_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[3] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[3]_i_1_n_0 ),
        .Q(\str_buffer_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[4] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[4]_i_1_n_0 ),
        .Q(p_1_in[0]));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[5] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[5]_i_1_n_0 ),
        .Q(p_1_in[1]));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[6] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[6]_i_1_n_0 ),
        .Q(p_0_in[0]));
  FDCE #(
    .INIT(1'b0)) 
    \str_buffer_reg[7] 
       (.C(md16_nd),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\str_buffer[7]_i_1_n_0 ),
        .Q(p_0_in[1]));
endmodule

(* ORIG_REF_NAME = "fifo4" *) 
module switch_elements_fifo4
   (DOB,
    E,
    D,
    clk_i,
    \wp_reg[0]_0 ,
    treg,
    out,
    \rp_reg[1]_0 ,
    \rp_reg[1]_1 ,
    Q,
    \dat_o_reg[7] ,
    wcol,
    spif,
    rst_i,
    \rp_reg[1]_2 ,
    \rp_reg[1]_3 ,
    \rp_reg[0]_0 );
  output [1:0]DOB;
  output [0:0]E;
  output [5:0]D;
  input clk_i;
  input \wp_reg[0]_0 ;
  input [7:0]treg;
  input out;
  input [1:0]\rp_reg[1]_0 ;
  input \rp_reg[1]_1 ;
  input [4:0]Q;
  input [5:0]\dat_o_reg[7] ;
  input wcol;
  input spif;
  input rst_i;
  input \rp_reg[1]_2 ;
  input \rp_reg[1]_3 ;
  input [0:0]\rp_reg[0]_0 ;

  wire [5:0]D;
  wire [1:0]DOB;
  wire [0:0]E;
  wire [4:0]Q;
  wire clk_i;
  wire [5:0]\dat_o_reg[7] ;
  wire [8:1]dout__0;
  wire gb;
  wire gb0;
  wire gb_i_1_n_0;
  wire out;
  wire p_14_in;
  wire rfempty;
  wire rffull;
  wire rfre;
  wire [1:0]rp;
  wire \rp[0]_i_1_n_0 ;
  wire \rp[1]_i_1_n_0 ;
  wire \rp[1]_i_2_n_0 ;
  wire [0:0]\rp_reg[0]_0 ;
  wire [1:0]\rp_reg[1]_0 ;
  wire \rp_reg[1]_1 ;
  wire \rp_reg[1]_2 ;
  wire \rp_reg[1]_3 ;
  wire rst_i;
  wire spif;
  wire [7:0]treg;
  wire wcol;
  wire [1:0]wp;
  wire \wp[0]_i_1_n_0 ;
  wire \wp[1]_i_2_n_0 ;
  wire \wp_reg[0]_0 ;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOE_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOF_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOG_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \dat_o[0]_i_1 
       (.I0(\dat_o_reg[7] [0]),
        .I1(rfempty),
        .I2(\rp_reg[1]_0 [0]),
        .I3(dout__0[1]),
        .I4(\rp_reg[1]_0 [1]),
        .I5(Q[0]),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'h00009009)) 
    \dat_o[0]_i_2 
       (.I0(rp[1]),
        .I1(wp[1]),
        .I2(rp[0]),
        .I3(wp[0]),
        .I4(gb),
        .O(rfempty));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \dat_o[1]_i_1 
       (.I0(\dat_o_reg[7] [1]),
        .I1(rffull),
        .I2(\rp_reg[1]_0 [0]),
        .I3(dout__0[2]),
        .I4(\rp_reg[1]_0 [1]),
        .I5(Q[1]),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'h90090000)) 
    \dat_o[1]_i_2 
       (.I0(rp[1]),
        .I1(wp[1]),
        .I2(rp[0]),
        .I3(wp[0]),
        .I4(gb),
        .O(rffull));
  LUT4 #(
    .INIT(16'hB833)) 
    \dat_o[4]_i_1 
       (.I0(\dat_o_reg[7] [2]),
        .I1(\rp_reg[1]_0 [0]),
        .I2(dout__0[5]),
        .I3(\rp_reg[1]_0 [1]),
        .O(D[2]));
  LUT5 #(
    .INIT(32'hB833B800)) 
    \dat_o[5]_i_1 
       (.I0(\dat_o_reg[7] [3]),
        .I1(\rp_reg[1]_0 [0]),
        .I2(dout__0[6]),
        .I3(\rp_reg[1]_0 [1]),
        .I4(Q[2]),
        .O(D[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \dat_o[6]_i_1 
       (.I0(\dat_o_reg[7] [4]),
        .I1(wcol),
        .I2(\rp_reg[1]_0 [0]),
        .I3(dout__0[7]),
        .I4(\rp_reg[1]_0 [1]),
        .I5(Q[3]),
        .O(D[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \dat_o[7]_i_1 
       (.I0(\dat_o_reg[7] [5]),
        .I1(spif),
        .I2(\rp_reg[1]_0 [0]),
        .I3(dout__0[8]),
        .I4(\rp_reg[1]_0 [1]),
        .I5(Q[4]),
        .O(D[5]));
  LUT5 #(
    .INIT(32'hF2000000)) 
    gb_i_1
       (.I0(gb),
        .I1(rfre),
        .I2(gb0),
        .I3(Q[3]),
        .I4(rst_i),
        .O(gb_i_1_n_0));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    gb_i_2__0
       (.I0(\rp_reg[1]_1 ),
        .I1(\rp_reg[1]_0 [0]),
        .I2(\rp_reg[1]_0 [1]),
        .I3(\rp_reg[1]_2 ),
        .I4(\rp_reg[1]_3 ),
        .I5(out),
        .O(rfre));
  LUT5 #(
    .INIT(32'h09600000)) 
    gb_i_3
       (.I0(rp[1]),
        .I1(wp[1]),
        .I2(wp[0]),
        .I3(rp[0]),
        .I4(\wp_reg[0]_0 ),
        .O(gb0));
  FDRE #(
    .INIT(1'b0)) 
    gb_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(gb_i_1_n_0),
        .Q(gb),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "32" *) 
  (* RTL_RAM_NAME = "rfifo/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "3" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "7" *) 
  RAM32M16_UNIQ_BASE_ mem_reg_0_3_0_7
       (.ADDRA({1'b0,1'b0,1'b0,rp}),
        .ADDRB({1'b0,1'b0,1'b0,rp}),
        .ADDRC({1'b0,1'b0,1'b0,rp}),
        .ADDRD({1'b0,1'b0,1'b0,rp}),
        .ADDRE({1'b0,1'b0,1'b0,rp}),
        .ADDRF({1'b0,1'b0,1'b0,rp}),
        .ADDRG({1'b0,1'b0,1'b0,rp}),
        .ADDRH({1'b0,1'b0,1'b0,wp}),
        .DIA(treg[1:0]),
        .DIB(treg[3:2]),
        .DIC(treg[5:4]),
        .DID(treg[7:6]),
        .DIE({1'b0,1'b0}),
        .DIF({1'b0,1'b0}),
        .DIG({1'b0,1'b0}),
        .DIH({1'b0,1'b0}),
        .DOA(dout__0[2:1]),
        .DOB(DOB),
        .DOC(dout__0[6:5]),
        .DOD(dout__0[8:7]),
        .DOE(NLW_mem_reg_0_3_0_7_DOE_UNCONNECTED[1:0]),
        .DOF(NLW_mem_reg_0_3_0_7_DOF_UNCONNECTED[1:0]),
        .DOG(NLW_mem_reg_0_3_0_7_DOG_UNCONNECTED[1:0]),
        .DOH(NLW_mem_reg_0_3_0_7_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(\wp_reg[0]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \rp[0]_i_1 
       (.I0(Q[3]),
        .I1(rp[0]),
        .O(\rp[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00400000FFFFFFFF)) 
    \rp[1]_i_1 
       (.I0(out),
        .I1(p_14_in),
        .I2(\rp_reg[1]_0 [1]),
        .I3(\rp_reg[1]_0 [0]),
        .I4(\rp_reg[1]_1 ),
        .I5(Q[3]),
        .O(\rp[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'h28)) 
    \rp[1]_i_2 
       (.I0(Q[3]),
        .I1(rp[1]),
        .I2(rp[0]),
        .O(\rp[1]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rp[1]_i_4 
       (.I0(\rp_reg[1]_2 ),
        .I1(\rp_reg[1]_3 ),
        .O(p_14_in));
  FDCE #(
    .INIT(1'b0)) 
    \rp_reg[0] 
       (.C(clk_i),
        .CE(\rp[1]_i_1_n_0 ),
        .CLR(\rp_reg[0]_0 ),
        .D(\rp[0]_i_1_n_0 ),
        .Q(rp[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rp_reg[1] 
       (.C(clk_i),
        .CE(\rp[1]_i_1_n_0 ),
        .CLR(\rp_reg[0]_0 ),
        .D(\rp[1]_i_2_n_0 ),
        .Q(rp[1]));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \wp[0]_i_1 
       (.I0(Q[3]),
        .I1(wp[0]),
        .O(\wp[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \wp[1]_i_1__0 
       (.I0(\wp_reg[0]_0 ),
        .I1(Q[3]),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \wp[1]_i_2 
       (.I0(wp[1]),
        .I1(wp[0]),
        .I2(Q[3]),
        .O(\wp[1]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \wp_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(\rp_reg[0]_0 ),
        .D(\wp[0]_i_1_n_0 ),
        .Q(wp[0]));
  FDCE #(
    .INIT(1'b0)) 
    \wp_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(\rp_reg[0]_0 ),
        .D(\wp[1]_i_2_n_0 ),
        .Q(wp[1]));
endmodule

(* ORIG_REF_NAME = "fifo4" *) 
module switch_elements_fifo4_5
   (\FSM_sequential_state_reg[1] ,
    \FSM_sequential_state_reg[0] ,
    D,
    \sper_reg[3] ,
    wcol0,
    E,
    clk_i,
    dat_i,
    sck_o_reg,
    Q,
    p_0_in,
    sck_o_reg_0,
    gb_reg_0,
    gb_reg_1,
    \treg_reg[7] ,
    \treg_reg[0] ,
    \dat_o_reg[3] ,
    \dat_o_reg[3]_0 ,
    DOB,
    rst_i,
    wcol,
    p_7_in,
    \wp_reg[1]_0 ,
    \wp_reg[1]_1 ,
    \wp_reg[1]_2 ,
    out,
    \wp_reg[0]_0 );
  output \FSM_sequential_state_reg[1] ;
  output \FSM_sequential_state_reg[0] ;
  output [7:0]D;
  output [1:0]\sper_reg[3] ;
  output wcol0;
  output [0:0]E;
  input clk_i;
  input [7:0]dat_i;
  input sck_o_reg;
  input [1:0]Q;
  input p_0_in;
  input sck_o_reg_0;
  input [2:0]gb_reg_0;
  input gb_reg_1;
  input [6:0]\treg_reg[7] ;
  input \treg_reg[0] ;
  input [1:0]\dat_o_reg[3] ;
  input [1:0]\dat_o_reg[3]_0 ;
  input [1:0]DOB;
  input rst_i;
  input wcol;
  input p_7_in;
  input \wp_reg[1]_0 ;
  input \wp_reg[1]_1 ;
  input \wp_reg[1]_2 ;
  input out;
  input [0:0]\wp_reg[0]_0 ;

  wire [7:0]D;
  wire [1:0]DOB;
  wire [0:0]E;
  wire \FSM_sequential_state_reg[0] ;
  wire \FSM_sequential_state_reg[1] ;
  wire [1:0]Q;
  wire clk_i;
  wire [7:0]dat_i;
  wire [1:0]\dat_o_reg[3] ;
  wire [1:0]\dat_o_reg[3]_0 ;
  wire [8:1]dout;
  wire gb;
  wire gb0;
  wire gb_i_1__0_n_0;
  wire [2:0]gb_reg_0;
  wire gb_reg_1;
  wire out;
  wire p_0_in;
  wire p_7_in;
  wire [1:0]rp;
  wire \rp[0]_i_1__0_n_0 ;
  wire \rp[1]_i_1__0_n_0 ;
  wire \rp[1]_i_2__0_n_0 ;
  wire rst_i;
  wire sck_o_i_2_n_0;
  wire sck_o_reg;
  wire sck_o_reg_0;
  wire [1:0]\sper_reg[3] ;
  wire \treg_reg[0] ;
  wire [6:0]\treg_reg[7] ;
  wire wcol;
  wire wcol0;
  wire wfempty;
  wire wffull;
  wire wfwe;
  wire [1:0]wp;
  wire \wp[0]_i_1__0_n_0 ;
  wire \wp[1]_i_1_n_0 ;
  wire \wp[1]_i_2__0_n_0 ;
  wire [0:0]\wp_reg[0]_0 ;
  wire \wp_reg[1]_0 ;
  wire \wp_reg[1]_1 ;
  wire \wp_reg[1]_2 ;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOE_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOF_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOG_UNCONNECTED;
  wire [1:0]NLW_mem_reg_0_3_0_7_DOH_UNCONNECTED;

  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'h0CC5)) 
    \FSM_sequential_state[1]_i_2 
       (.I0(wfempty),
        .I1(p_0_in),
        .I2(Q[0]),
        .I3(Q[1]),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'h00009009)) 
    \FSM_sequential_state[1]_i_4 
       (.I0(rp[1]),
        .I1(wp[1]),
        .I2(rp[0]),
        .I3(wp[0]),
        .I4(gb),
        .O(wfempty));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \dat_o[2]_i_1 
       (.I0(\dat_o_reg[3] [0]),
        .I1(wfempty),
        .I2(\dat_o_reg[3]_0 [0]),
        .I3(DOB[0]),
        .I4(\dat_o_reg[3]_0 [1]),
        .I5(gb_reg_0[0]),
        .O(\sper_reg[3] [0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \dat_o[3]_i_1 
       (.I0(\dat_o_reg[3] [1]),
        .I1(wffull),
        .I2(\dat_o_reg[3]_0 [0]),
        .I3(DOB[1]),
        .I4(\dat_o_reg[3]_0 [1]),
        .I5(gb_reg_0[1]),
        .O(\sper_reg[3] [1]));
  LUT5 #(
    .INIT(32'hF2000000)) 
    gb_i_1__0
       (.I0(gb),
        .I1(gb_reg_1),
        .I2(gb0),
        .I3(gb_reg_0[2]),
        .I4(rst_i),
        .O(gb_i_1__0_n_0));
  LUT5 #(
    .INIT(32'h09600000)) 
    gb_i_2
       (.I0(rp[1]),
        .I1(wp[1]),
        .I2(wp[0]),
        .I3(rp[0]),
        .I4(wfwe),
        .O(gb0));
  FDRE #(
    .INIT(1'b0)) 
    gb_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(gb_i_1__0_n_0),
        .Q(gb),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "32" *) 
  (* RTL_RAM_NAME = "wfifo/mem" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "3" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "7" *) 
  RAM32M16_HD32711 mem_reg_0_3_0_7
       (.ADDRA({1'b0,1'b0,1'b0,rp}),
        .ADDRB({1'b0,1'b0,1'b0,rp}),
        .ADDRC({1'b0,1'b0,1'b0,rp}),
        .ADDRD({1'b0,1'b0,1'b0,rp}),
        .ADDRE({1'b0,1'b0,1'b0,rp}),
        .ADDRF({1'b0,1'b0,1'b0,rp}),
        .ADDRG({1'b0,1'b0,1'b0,rp}),
        .ADDRH({1'b0,1'b0,1'b0,wp}),
        .DIA(dat_i[1:0]),
        .DIB(dat_i[3:2]),
        .DIC(dat_i[5:4]),
        .DID(dat_i[7:6]),
        .DIE({1'b0,1'b0}),
        .DIF({1'b0,1'b0}),
        .DIG({1'b0,1'b0}),
        .DIH({1'b0,1'b0}),
        .DOA(dout[2:1]),
        .DOB(dout[4:3]),
        .DOC(dout[6:5]),
        .DOD(dout[8:7]),
        .DOE(NLW_mem_reg_0_3_0_7_DOE_UNCONNECTED[1:0]),
        .DOF(NLW_mem_reg_0_3_0_7_DOF_UNCONNECTED[1:0]),
        .DOG(NLW_mem_reg_0_3_0_7_DOG_UNCONNECTED[1:0]),
        .DOH(NLW_mem_reg_0_3_0_7_DOH_UNCONNECTED[1:0]),
        .WCLK(clk_i),
        .WE(wfwe));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    mem_reg_0_3_0_7_i_1
       (.I0(\wp_reg[1]_0 ),
        .I1(\dat_o_reg[3]_0 [0]),
        .I2(\dat_o_reg[3]_0 [1]),
        .I3(\wp_reg[1]_1 ),
        .I4(\wp_reg[1]_2 ),
        .I5(out),
        .O(wfwe));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \rp[0]_i_1__0 
       (.I0(gb_reg_0[2]),
        .I1(rp[0]),
        .O(\rp[0]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rp[1]_i_1__0 
       (.I0(gb_reg_1),
        .I1(gb_reg_0[2]),
        .O(\rp[1]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'h28)) 
    \rp[1]_i_2__0 
       (.I0(gb_reg_0[2]),
        .I1(rp[1]),
        .I2(rp[0]),
        .O(\rp[1]_i_2__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \rp_reg[0] 
       (.C(clk_i),
        .CE(\rp[1]_i_1__0_n_0 ),
        .CLR(\wp_reg[0]_0 ),
        .D(\rp[0]_i_1__0_n_0 ),
        .Q(rp[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rp_reg[1] 
       (.C(clk_i),
        .CE(\rp[1]_i_1__0_n_0 ),
        .CLR(\wp_reg[0]_0 ),
        .D(\rp[1]_i_2__0_n_0 ),
        .Q(rp[1]));
  LUT6 #(
    .INIT(64'hFAFFEAFA0F00EA0A)) 
    sck_o_i_1
       (.I0(sck_o_i_2_n_0),
        .I1(sck_o_reg),
        .I2(Q[1]),
        .I3(p_0_in),
        .I4(Q[0]),
        .I5(sck_o_reg_0),
        .O(\FSM_sequential_state_reg[1] ));
  LUT6 #(
    .INIT(64'h000000000000AA2E)) 
    sck_o_i_2
       (.I0(gb_reg_0[1]),
        .I1(gb_reg_0[0]),
        .I2(sck_o_reg_0),
        .I3(wfempty),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(sck_o_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[0]_i_1 
       (.I0(dout[1]),
        .I1(Q[1]),
        .I2(\treg_reg[0] ),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[1]_i_1 
       (.I0(dout[2]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [0]),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[2]_i_1 
       (.I0(dout[3]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [1]),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[3]_i_1 
       (.I0(dout[4]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [2]),
        .O(D[3]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[4]_i_1 
       (.I0(dout[5]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [3]),
        .O(D[4]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[5]_i_1 
       (.I0(dout[6]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [4]),
        .O(D[5]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[6]_i_1 
       (.I0(dout[7]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [5]),
        .O(D[6]));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \treg[7]_i_2 
       (.I0(dout[8]),
        .I1(Q[1]),
        .I2(\treg_reg[7] [6]),
        .O(D[7]));
  LUT5 #(
    .INIT(32'h00EAEAEA)) 
    wcol_i_1
       (.I0(wcol),
        .I1(wfwe),
        .I2(wffull),
        .I3(dat_i[6]),
        .I4(p_7_in),
        .O(wcol0));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'h90090000)) 
    wcol_i_2
       (.I0(rp[1]),
        .I1(wp[1]),
        .I2(rp[0]),
        .I3(wp[0]),
        .I4(gb),
        .O(wffull));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'h01)) 
    wfre_i_1
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(wfempty),
        .O(\FSM_sequential_state_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \wp[0]_i_1__0 
       (.I0(gb_reg_0[2]),
        .I1(wp[0]),
        .O(\wp[0]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \wp[1]_i_1 
       (.I0(wfwe),
        .I1(gb_reg_0[2]),
        .O(\wp[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \wp[1]_i_2__0 
       (.I0(wp[1]),
        .I1(wp[0]),
        .I2(gb_reg_0[2]),
        .O(\wp[1]_i_2__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \wp_reg[0] 
       (.C(clk_i),
        .CE(\wp[1]_i_1_n_0 ),
        .CLR(\wp_reg[0]_0 ),
        .D(\wp[0]_i_1__0_n_0 ),
        .Q(wp[0]));
  FDCE #(
    .INIT(1'b0)) 
    \wp_reg[1] 
       (.C(clk_i),
        .CE(\wp[1]_i_1_n_0 ),
        .CLR(\wp_reg[0]_0 ),
        .D(\wp[1]_i_2__0_n_0 ),
        .Q(wp[1]));
endmodule

(* ORIG_REF_NAME = "manage_registers" *) 
module switch_elements_manage_registers
   (in0,
    mdio_out_valid,
    Q,
    cfgRxRegData,
    cfgTxRegData,
    mgmt_rd_data,
    mdio_opcode,
    mdio_in_valid,
    clk_i,
    rst_i,
    out,
    \stat_rd_data_reg[63]_0 ,
    \stat_rd_data_reg[63]_1 ,
    \recv_config0_reg[0]_0 ,
    \mgmt_rd_data_reg[15]_0 ,
    mgmt_wr_data,
    rxStatRegPlus,
    txStatRegPlus);
  output in0;
  output mdio_out_valid;
  output [4:0]Q;
  output [52:0]cfgRxRegData;
  output [9:0]cfgTxRegData;
  output [31:0]mgmt_rd_data;
  output [0:0]mdio_opcode;
  input mdio_in_valid;
  input clk_i;
  input rst_i;
  input [9:0]out;
  input \stat_rd_data_reg[63]_0 ;
  input \stat_rd_data_reg[63]_1 ;
  input [0:0]\recv_config0_reg[0]_0 ;
  input [15:0]\mgmt_rd_data_reg[15]_0 ;
  input [31:0]mgmt_wr_data;
  input [18:0]rxStatRegPlus;
  input [14:0]txStatRegPlus;

  wire [4:0]Q;
  wire \broadcast_frame_transed[0]_i_2_n_0 ;
  wire [63:0]broadcast_frame_transed_reg;
  wire \broadcast_frame_transed_reg[0]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[0]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[16]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[24]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[32]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[40]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[48]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[56]_i_1_n_9 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_0 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_1 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_10 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_11 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_12 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_13 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_14 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_15 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_2 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_3 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_4 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_5 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_6 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_7 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_8 ;
  wire \broadcast_frame_transed_reg[8]_i_1_n_9 ;
  wire \broadcast_received_good[0]_i_2_n_0 ;
  wire [63:0]broadcast_received_good_reg;
  wire \broadcast_received_good_reg[0]_i_1_n_0 ;
  wire \broadcast_received_good_reg[0]_i_1_n_1 ;
  wire \broadcast_received_good_reg[0]_i_1_n_10 ;
  wire \broadcast_received_good_reg[0]_i_1_n_11 ;
  wire \broadcast_received_good_reg[0]_i_1_n_12 ;
  wire \broadcast_received_good_reg[0]_i_1_n_13 ;
  wire \broadcast_received_good_reg[0]_i_1_n_14 ;
  wire \broadcast_received_good_reg[0]_i_1_n_15 ;
  wire \broadcast_received_good_reg[0]_i_1_n_2 ;
  wire \broadcast_received_good_reg[0]_i_1_n_3 ;
  wire \broadcast_received_good_reg[0]_i_1_n_4 ;
  wire \broadcast_received_good_reg[0]_i_1_n_5 ;
  wire \broadcast_received_good_reg[0]_i_1_n_6 ;
  wire \broadcast_received_good_reg[0]_i_1_n_7 ;
  wire \broadcast_received_good_reg[0]_i_1_n_8 ;
  wire \broadcast_received_good_reg[0]_i_1_n_9 ;
  wire \broadcast_received_good_reg[16]_i_1_n_0 ;
  wire \broadcast_received_good_reg[16]_i_1_n_1 ;
  wire \broadcast_received_good_reg[16]_i_1_n_10 ;
  wire \broadcast_received_good_reg[16]_i_1_n_11 ;
  wire \broadcast_received_good_reg[16]_i_1_n_12 ;
  wire \broadcast_received_good_reg[16]_i_1_n_13 ;
  wire \broadcast_received_good_reg[16]_i_1_n_14 ;
  wire \broadcast_received_good_reg[16]_i_1_n_15 ;
  wire \broadcast_received_good_reg[16]_i_1_n_2 ;
  wire \broadcast_received_good_reg[16]_i_1_n_3 ;
  wire \broadcast_received_good_reg[16]_i_1_n_4 ;
  wire \broadcast_received_good_reg[16]_i_1_n_5 ;
  wire \broadcast_received_good_reg[16]_i_1_n_6 ;
  wire \broadcast_received_good_reg[16]_i_1_n_7 ;
  wire \broadcast_received_good_reg[16]_i_1_n_8 ;
  wire \broadcast_received_good_reg[16]_i_1_n_9 ;
  wire \broadcast_received_good_reg[24]_i_1_n_0 ;
  wire \broadcast_received_good_reg[24]_i_1_n_1 ;
  wire \broadcast_received_good_reg[24]_i_1_n_10 ;
  wire \broadcast_received_good_reg[24]_i_1_n_11 ;
  wire \broadcast_received_good_reg[24]_i_1_n_12 ;
  wire \broadcast_received_good_reg[24]_i_1_n_13 ;
  wire \broadcast_received_good_reg[24]_i_1_n_14 ;
  wire \broadcast_received_good_reg[24]_i_1_n_15 ;
  wire \broadcast_received_good_reg[24]_i_1_n_2 ;
  wire \broadcast_received_good_reg[24]_i_1_n_3 ;
  wire \broadcast_received_good_reg[24]_i_1_n_4 ;
  wire \broadcast_received_good_reg[24]_i_1_n_5 ;
  wire \broadcast_received_good_reg[24]_i_1_n_6 ;
  wire \broadcast_received_good_reg[24]_i_1_n_7 ;
  wire \broadcast_received_good_reg[24]_i_1_n_8 ;
  wire \broadcast_received_good_reg[24]_i_1_n_9 ;
  wire \broadcast_received_good_reg[32]_i_1_n_0 ;
  wire \broadcast_received_good_reg[32]_i_1_n_1 ;
  wire \broadcast_received_good_reg[32]_i_1_n_10 ;
  wire \broadcast_received_good_reg[32]_i_1_n_11 ;
  wire \broadcast_received_good_reg[32]_i_1_n_12 ;
  wire \broadcast_received_good_reg[32]_i_1_n_13 ;
  wire \broadcast_received_good_reg[32]_i_1_n_14 ;
  wire \broadcast_received_good_reg[32]_i_1_n_15 ;
  wire \broadcast_received_good_reg[32]_i_1_n_2 ;
  wire \broadcast_received_good_reg[32]_i_1_n_3 ;
  wire \broadcast_received_good_reg[32]_i_1_n_4 ;
  wire \broadcast_received_good_reg[32]_i_1_n_5 ;
  wire \broadcast_received_good_reg[32]_i_1_n_6 ;
  wire \broadcast_received_good_reg[32]_i_1_n_7 ;
  wire \broadcast_received_good_reg[32]_i_1_n_8 ;
  wire \broadcast_received_good_reg[32]_i_1_n_9 ;
  wire \broadcast_received_good_reg[40]_i_1_n_0 ;
  wire \broadcast_received_good_reg[40]_i_1_n_1 ;
  wire \broadcast_received_good_reg[40]_i_1_n_10 ;
  wire \broadcast_received_good_reg[40]_i_1_n_11 ;
  wire \broadcast_received_good_reg[40]_i_1_n_12 ;
  wire \broadcast_received_good_reg[40]_i_1_n_13 ;
  wire \broadcast_received_good_reg[40]_i_1_n_14 ;
  wire \broadcast_received_good_reg[40]_i_1_n_15 ;
  wire \broadcast_received_good_reg[40]_i_1_n_2 ;
  wire \broadcast_received_good_reg[40]_i_1_n_3 ;
  wire \broadcast_received_good_reg[40]_i_1_n_4 ;
  wire \broadcast_received_good_reg[40]_i_1_n_5 ;
  wire \broadcast_received_good_reg[40]_i_1_n_6 ;
  wire \broadcast_received_good_reg[40]_i_1_n_7 ;
  wire \broadcast_received_good_reg[40]_i_1_n_8 ;
  wire \broadcast_received_good_reg[40]_i_1_n_9 ;
  wire \broadcast_received_good_reg[48]_i_1_n_0 ;
  wire \broadcast_received_good_reg[48]_i_1_n_1 ;
  wire \broadcast_received_good_reg[48]_i_1_n_10 ;
  wire \broadcast_received_good_reg[48]_i_1_n_11 ;
  wire \broadcast_received_good_reg[48]_i_1_n_12 ;
  wire \broadcast_received_good_reg[48]_i_1_n_13 ;
  wire \broadcast_received_good_reg[48]_i_1_n_14 ;
  wire \broadcast_received_good_reg[48]_i_1_n_15 ;
  wire \broadcast_received_good_reg[48]_i_1_n_2 ;
  wire \broadcast_received_good_reg[48]_i_1_n_3 ;
  wire \broadcast_received_good_reg[48]_i_1_n_4 ;
  wire \broadcast_received_good_reg[48]_i_1_n_5 ;
  wire \broadcast_received_good_reg[48]_i_1_n_6 ;
  wire \broadcast_received_good_reg[48]_i_1_n_7 ;
  wire \broadcast_received_good_reg[48]_i_1_n_8 ;
  wire \broadcast_received_good_reg[48]_i_1_n_9 ;
  wire \broadcast_received_good_reg[56]_i_1_n_1 ;
  wire \broadcast_received_good_reg[56]_i_1_n_10 ;
  wire \broadcast_received_good_reg[56]_i_1_n_11 ;
  wire \broadcast_received_good_reg[56]_i_1_n_12 ;
  wire \broadcast_received_good_reg[56]_i_1_n_13 ;
  wire \broadcast_received_good_reg[56]_i_1_n_14 ;
  wire \broadcast_received_good_reg[56]_i_1_n_15 ;
  wire \broadcast_received_good_reg[56]_i_1_n_2 ;
  wire \broadcast_received_good_reg[56]_i_1_n_3 ;
  wire \broadcast_received_good_reg[56]_i_1_n_4 ;
  wire \broadcast_received_good_reg[56]_i_1_n_5 ;
  wire \broadcast_received_good_reg[56]_i_1_n_6 ;
  wire \broadcast_received_good_reg[56]_i_1_n_7 ;
  wire \broadcast_received_good_reg[56]_i_1_n_8 ;
  wire \broadcast_received_good_reg[56]_i_1_n_9 ;
  wire \broadcast_received_good_reg[8]_i_1_n_0 ;
  wire \broadcast_received_good_reg[8]_i_1_n_1 ;
  wire \broadcast_received_good_reg[8]_i_1_n_10 ;
  wire \broadcast_received_good_reg[8]_i_1_n_11 ;
  wire \broadcast_received_good_reg[8]_i_1_n_12 ;
  wire \broadcast_received_good_reg[8]_i_1_n_13 ;
  wire \broadcast_received_good_reg[8]_i_1_n_14 ;
  wire \broadcast_received_good_reg[8]_i_1_n_15 ;
  wire \broadcast_received_good_reg[8]_i_1_n_2 ;
  wire \broadcast_received_good_reg[8]_i_1_n_3 ;
  wire \broadcast_received_good_reg[8]_i_1_n_4 ;
  wire \broadcast_received_good_reg[8]_i_1_n_5 ;
  wire \broadcast_received_good_reg[8]_i_1_n_6 ;
  wire \broadcast_received_good_reg[8]_i_1_n_7 ;
  wire \broadcast_received_good_reg[8]_i_1_n_8 ;
  wire \broadcast_received_good_reg[8]_i_1_n_9 ;
  wire [52:0]cfgRxRegData;
  wire [9:0]cfgTxRegData;
  wire clk_i;
  wire \control_frame_good[0]_i_2_n_0 ;
  wire [63:0]control_frame_good_reg;
  wire \control_frame_good_reg[0]_i_1_n_0 ;
  wire \control_frame_good_reg[0]_i_1_n_1 ;
  wire \control_frame_good_reg[0]_i_1_n_10 ;
  wire \control_frame_good_reg[0]_i_1_n_11 ;
  wire \control_frame_good_reg[0]_i_1_n_12 ;
  wire \control_frame_good_reg[0]_i_1_n_13 ;
  wire \control_frame_good_reg[0]_i_1_n_14 ;
  wire \control_frame_good_reg[0]_i_1_n_15 ;
  wire \control_frame_good_reg[0]_i_1_n_2 ;
  wire \control_frame_good_reg[0]_i_1_n_3 ;
  wire \control_frame_good_reg[0]_i_1_n_4 ;
  wire \control_frame_good_reg[0]_i_1_n_5 ;
  wire \control_frame_good_reg[0]_i_1_n_6 ;
  wire \control_frame_good_reg[0]_i_1_n_7 ;
  wire \control_frame_good_reg[0]_i_1_n_8 ;
  wire \control_frame_good_reg[0]_i_1_n_9 ;
  wire \control_frame_good_reg[16]_i_1_n_0 ;
  wire \control_frame_good_reg[16]_i_1_n_1 ;
  wire \control_frame_good_reg[16]_i_1_n_10 ;
  wire \control_frame_good_reg[16]_i_1_n_11 ;
  wire \control_frame_good_reg[16]_i_1_n_12 ;
  wire \control_frame_good_reg[16]_i_1_n_13 ;
  wire \control_frame_good_reg[16]_i_1_n_14 ;
  wire \control_frame_good_reg[16]_i_1_n_15 ;
  wire \control_frame_good_reg[16]_i_1_n_2 ;
  wire \control_frame_good_reg[16]_i_1_n_3 ;
  wire \control_frame_good_reg[16]_i_1_n_4 ;
  wire \control_frame_good_reg[16]_i_1_n_5 ;
  wire \control_frame_good_reg[16]_i_1_n_6 ;
  wire \control_frame_good_reg[16]_i_1_n_7 ;
  wire \control_frame_good_reg[16]_i_1_n_8 ;
  wire \control_frame_good_reg[16]_i_1_n_9 ;
  wire \control_frame_good_reg[24]_i_1_n_0 ;
  wire \control_frame_good_reg[24]_i_1_n_1 ;
  wire \control_frame_good_reg[24]_i_1_n_10 ;
  wire \control_frame_good_reg[24]_i_1_n_11 ;
  wire \control_frame_good_reg[24]_i_1_n_12 ;
  wire \control_frame_good_reg[24]_i_1_n_13 ;
  wire \control_frame_good_reg[24]_i_1_n_14 ;
  wire \control_frame_good_reg[24]_i_1_n_15 ;
  wire \control_frame_good_reg[24]_i_1_n_2 ;
  wire \control_frame_good_reg[24]_i_1_n_3 ;
  wire \control_frame_good_reg[24]_i_1_n_4 ;
  wire \control_frame_good_reg[24]_i_1_n_5 ;
  wire \control_frame_good_reg[24]_i_1_n_6 ;
  wire \control_frame_good_reg[24]_i_1_n_7 ;
  wire \control_frame_good_reg[24]_i_1_n_8 ;
  wire \control_frame_good_reg[24]_i_1_n_9 ;
  wire \control_frame_good_reg[32]_i_1_n_0 ;
  wire \control_frame_good_reg[32]_i_1_n_1 ;
  wire \control_frame_good_reg[32]_i_1_n_10 ;
  wire \control_frame_good_reg[32]_i_1_n_11 ;
  wire \control_frame_good_reg[32]_i_1_n_12 ;
  wire \control_frame_good_reg[32]_i_1_n_13 ;
  wire \control_frame_good_reg[32]_i_1_n_14 ;
  wire \control_frame_good_reg[32]_i_1_n_15 ;
  wire \control_frame_good_reg[32]_i_1_n_2 ;
  wire \control_frame_good_reg[32]_i_1_n_3 ;
  wire \control_frame_good_reg[32]_i_1_n_4 ;
  wire \control_frame_good_reg[32]_i_1_n_5 ;
  wire \control_frame_good_reg[32]_i_1_n_6 ;
  wire \control_frame_good_reg[32]_i_1_n_7 ;
  wire \control_frame_good_reg[32]_i_1_n_8 ;
  wire \control_frame_good_reg[32]_i_1_n_9 ;
  wire \control_frame_good_reg[40]_i_1_n_0 ;
  wire \control_frame_good_reg[40]_i_1_n_1 ;
  wire \control_frame_good_reg[40]_i_1_n_10 ;
  wire \control_frame_good_reg[40]_i_1_n_11 ;
  wire \control_frame_good_reg[40]_i_1_n_12 ;
  wire \control_frame_good_reg[40]_i_1_n_13 ;
  wire \control_frame_good_reg[40]_i_1_n_14 ;
  wire \control_frame_good_reg[40]_i_1_n_15 ;
  wire \control_frame_good_reg[40]_i_1_n_2 ;
  wire \control_frame_good_reg[40]_i_1_n_3 ;
  wire \control_frame_good_reg[40]_i_1_n_4 ;
  wire \control_frame_good_reg[40]_i_1_n_5 ;
  wire \control_frame_good_reg[40]_i_1_n_6 ;
  wire \control_frame_good_reg[40]_i_1_n_7 ;
  wire \control_frame_good_reg[40]_i_1_n_8 ;
  wire \control_frame_good_reg[40]_i_1_n_9 ;
  wire \control_frame_good_reg[48]_i_1_n_0 ;
  wire \control_frame_good_reg[48]_i_1_n_1 ;
  wire \control_frame_good_reg[48]_i_1_n_10 ;
  wire \control_frame_good_reg[48]_i_1_n_11 ;
  wire \control_frame_good_reg[48]_i_1_n_12 ;
  wire \control_frame_good_reg[48]_i_1_n_13 ;
  wire \control_frame_good_reg[48]_i_1_n_14 ;
  wire \control_frame_good_reg[48]_i_1_n_15 ;
  wire \control_frame_good_reg[48]_i_1_n_2 ;
  wire \control_frame_good_reg[48]_i_1_n_3 ;
  wire \control_frame_good_reg[48]_i_1_n_4 ;
  wire \control_frame_good_reg[48]_i_1_n_5 ;
  wire \control_frame_good_reg[48]_i_1_n_6 ;
  wire \control_frame_good_reg[48]_i_1_n_7 ;
  wire \control_frame_good_reg[48]_i_1_n_8 ;
  wire \control_frame_good_reg[48]_i_1_n_9 ;
  wire \control_frame_good_reg[56]_i_1_n_1 ;
  wire \control_frame_good_reg[56]_i_1_n_10 ;
  wire \control_frame_good_reg[56]_i_1_n_11 ;
  wire \control_frame_good_reg[56]_i_1_n_12 ;
  wire \control_frame_good_reg[56]_i_1_n_13 ;
  wire \control_frame_good_reg[56]_i_1_n_14 ;
  wire \control_frame_good_reg[56]_i_1_n_15 ;
  wire \control_frame_good_reg[56]_i_1_n_2 ;
  wire \control_frame_good_reg[56]_i_1_n_3 ;
  wire \control_frame_good_reg[56]_i_1_n_4 ;
  wire \control_frame_good_reg[56]_i_1_n_5 ;
  wire \control_frame_good_reg[56]_i_1_n_6 ;
  wire \control_frame_good_reg[56]_i_1_n_7 ;
  wire \control_frame_good_reg[56]_i_1_n_8 ;
  wire \control_frame_good_reg[56]_i_1_n_9 ;
  wire \control_frame_good_reg[8]_i_1_n_0 ;
  wire \control_frame_good_reg[8]_i_1_n_1 ;
  wire \control_frame_good_reg[8]_i_1_n_10 ;
  wire \control_frame_good_reg[8]_i_1_n_11 ;
  wire \control_frame_good_reg[8]_i_1_n_12 ;
  wire \control_frame_good_reg[8]_i_1_n_13 ;
  wire \control_frame_good_reg[8]_i_1_n_14 ;
  wire \control_frame_good_reg[8]_i_1_n_15 ;
  wire \control_frame_good_reg[8]_i_1_n_2 ;
  wire \control_frame_good_reg[8]_i_1_n_3 ;
  wire \control_frame_good_reg[8]_i_1_n_4 ;
  wire \control_frame_good_reg[8]_i_1_n_5 ;
  wire \control_frame_good_reg[8]_i_1_n_6 ;
  wire \control_frame_good_reg[8]_i_1_n_7 ;
  wire \control_frame_good_reg[8]_i_1_n_8 ;
  wire \control_frame_good_reg[8]_i_1_n_9 ;
  wire \control_frame_transed[0]_i_2_n_0 ;
  wire [63:0]control_frame_transed_reg;
  wire \control_frame_transed_reg[0]_i_1_n_0 ;
  wire \control_frame_transed_reg[0]_i_1_n_1 ;
  wire \control_frame_transed_reg[0]_i_1_n_10 ;
  wire \control_frame_transed_reg[0]_i_1_n_11 ;
  wire \control_frame_transed_reg[0]_i_1_n_12 ;
  wire \control_frame_transed_reg[0]_i_1_n_13 ;
  wire \control_frame_transed_reg[0]_i_1_n_14 ;
  wire \control_frame_transed_reg[0]_i_1_n_15 ;
  wire \control_frame_transed_reg[0]_i_1_n_2 ;
  wire \control_frame_transed_reg[0]_i_1_n_3 ;
  wire \control_frame_transed_reg[0]_i_1_n_4 ;
  wire \control_frame_transed_reg[0]_i_1_n_5 ;
  wire \control_frame_transed_reg[0]_i_1_n_6 ;
  wire \control_frame_transed_reg[0]_i_1_n_7 ;
  wire \control_frame_transed_reg[0]_i_1_n_8 ;
  wire \control_frame_transed_reg[0]_i_1_n_9 ;
  wire \control_frame_transed_reg[16]_i_1_n_0 ;
  wire \control_frame_transed_reg[16]_i_1_n_1 ;
  wire \control_frame_transed_reg[16]_i_1_n_10 ;
  wire \control_frame_transed_reg[16]_i_1_n_11 ;
  wire \control_frame_transed_reg[16]_i_1_n_12 ;
  wire \control_frame_transed_reg[16]_i_1_n_13 ;
  wire \control_frame_transed_reg[16]_i_1_n_14 ;
  wire \control_frame_transed_reg[16]_i_1_n_15 ;
  wire \control_frame_transed_reg[16]_i_1_n_2 ;
  wire \control_frame_transed_reg[16]_i_1_n_3 ;
  wire \control_frame_transed_reg[16]_i_1_n_4 ;
  wire \control_frame_transed_reg[16]_i_1_n_5 ;
  wire \control_frame_transed_reg[16]_i_1_n_6 ;
  wire \control_frame_transed_reg[16]_i_1_n_7 ;
  wire \control_frame_transed_reg[16]_i_1_n_8 ;
  wire \control_frame_transed_reg[16]_i_1_n_9 ;
  wire \control_frame_transed_reg[24]_i_1_n_0 ;
  wire \control_frame_transed_reg[24]_i_1_n_1 ;
  wire \control_frame_transed_reg[24]_i_1_n_10 ;
  wire \control_frame_transed_reg[24]_i_1_n_11 ;
  wire \control_frame_transed_reg[24]_i_1_n_12 ;
  wire \control_frame_transed_reg[24]_i_1_n_13 ;
  wire \control_frame_transed_reg[24]_i_1_n_14 ;
  wire \control_frame_transed_reg[24]_i_1_n_15 ;
  wire \control_frame_transed_reg[24]_i_1_n_2 ;
  wire \control_frame_transed_reg[24]_i_1_n_3 ;
  wire \control_frame_transed_reg[24]_i_1_n_4 ;
  wire \control_frame_transed_reg[24]_i_1_n_5 ;
  wire \control_frame_transed_reg[24]_i_1_n_6 ;
  wire \control_frame_transed_reg[24]_i_1_n_7 ;
  wire \control_frame_transed_reg[24]_i_1_n_8 ;
  wire \control_frame_transed_reg[24]_i_1_n_9 ;
  wire \control_frame_transed_reg[32]_i_1_n_0 ;
  wire \control_frame_transed_reg[32]_i_1_n_1 ;
  wire \control_frame_transed_reg[32]_i_1_n_10 ;
  wire \control_frame_transed_reg[32]_i_1_n_11 ;
  wire \control_frame_transed_reg[32]_i_1_n_12 ;
  wire \control_frame_transed_reg[32]_i_1_n_13 ;
  wire \control_frame_transed_reg[32]_i_1_n_14 ;
  wire \control_frame_transed_reg[32]_i_1_n_15 ;
  wire \control_frame_transed_reg[32]_i_1_n_2 ;
  wire \control_frame_transed_reg[32]_i_1_n_3 ;
  wire \control_frame_transed_reg[32]_i_1_n_4 ;
  wire \control_frame_transed_reg[32]_i_1_n_5 ;
  wire \control_frame_transed_reg[32]_i_1_n_6 ;
  wire \control_frame_transed_reg[32]_i_1_n_7 ;
  wire \control_frame_transed_reg[32]_i_1_n_8 ;
  wire \control_frame_transed_reg[32]_i_1_n_9 ;
  wire \control_frame_transed_reg[40]_i_1_n_0 ;
  wire \control_frame_transed_reg[40]_i_1_n_1 ;
  wire \control_frame_transed_reg[40]_i_1_n_10 ;
  wire \control_frame_transed_reg[40]_i_1_n_11 ;
  wire \control_frame_transed_reg[40]_i_1_n_12 ;
  wire \control_frame_transed_reg[40]_i_1_n_13 ;
  wire \control_frame_transed_reg[40]_i_1_n_14 ;
  wire \control_frame_transed_reg[40]_i_1_n_15 ;
  wire \control_frame_transed_reg[40]_i_1_n_2 ;
  wire \control_frame_transed_reg[40]_i_1_n_3 ;
  wire \control_frame_transed_reg[40]_i_1_n_4 ;
  wire \control_frame_transed_reg[40]_i_1_n_5 ;
  wire \control_frame_transed_reg[40]_i_1_n_6 ;
  wire \control_frame_transed_reg[40]_i_1_n_7 ;
  wire \control_frame_transed_reg[40]_i_1_n_8 ;
  wire \control_frame_transed_reg[40]_i_1_n_9 ;
  wire \control_frame_transed_reg[48]_i_1_n_0 ;
  wire \control_frame_transed_reg[48]_i_1_n_1 ;
  wire \control_frame_transed_reg[48]_i_1_n_10 ;
  wire \control_frame_transed_reg[48]_i_1_n_11 ;
  wire \control_frame_transed_reg[48]_i_1_n_12 ;
  wire \control_frame_transed_reg[48]_i_1_n_13 ;
  wire \control_frame_transed_reg[48]_i_1_n_14 ;
  wire \control_frame_transed_reg[48]_i_1_n_15 ;
  wire \control_frame_transed_reg[48]_i_1_n_2 ;
  wire \control_frame_transed_reg[48]_i_1_n_3 ;
  wire \control_frame_transed_reg[48]_i_1_n_4 ;
  wire \control_frame_transed_reg[48]_i_1_n_5 ;
  wire \control_frame_transed_reg[48]_i_1_n_6 ;
  wire \control_frame_transed_reg[48]_i_1_n_7 ;
  wire \control_frame_transed_reg[48]_i_1_n_8 ;
  wire \control_frame_transed_reg[48]_i_1_n_9 ;
  wire \control_frame_transed_reg[56]_i_1_n_1 ;
  wire \control_frame_transed_reg[56]_i_1_n_10 ;
  wire \control_frame_transed_reg[56]_i_1_n_11 ;
  wire \control_frame_transed_reg[56]_i_1_n_12 ;
  wire \control_frame_transed_reg[56]_i_1_n_13 ;
  wire \control_frame_transed_reg[56]_i_1_n_14 ;
  wire \control_frame_transed_reg[56]_i_1_n_15 ;
  wire \control_frame_transed_reg[56]_i_1_n_2 ;
  wire \control_frame_transed_reg[56]_i_1_n_3 ;
  wire \control_frame_transed_reg[56]_i_1_n_4 ;
  wire \control_frame_transed_reg[56]_i_1_n_5 ;
  wire \control_frame_transed_reg[56]_i_1_n_6 ;
  wire \control_frame_transed_reg[56]_i_1_n_7 ;
  wire \control_frame_transed_reg[56]_i_1_n_8 ;
  wire \control_frame_transed_reg[56]_i_1_n_9 ;
  wire \control_frame_transed_reg[8]_i_1_n_0 ;
  wire \control_frame_transed_reg[8]_i_1_n_1 ;
  wire \control_frame_transed_reg[8]_i_1_n_10 ;
  wire \control_frame_transed_reg[8]_i_1_n_11 ;
  wire \control_frame_transed_reg[8]_i_1_n_12 ;
  wire \control_frame_transed_reg[8]_i_1_n_13 ;
  wire \control_frame_transed_reg[8]_i_1_n_14 ;
  wire \control_frame_transed_reg[8]_i_1_n_15 ;
  wire \control_frame_transed_reg[8]_i_1_n_2 ;
  wire \control_frame_transed_reg[8]_i_1_n_3 ;
  wire \control_frame_transed_reg[8]_i_1_n_4 ;
  wire \control_frame_transed_reg[8]_i_1_n_5 ;
  wire \control_frame_transed_reg[8]_i_1_n_6 ;
  wire \control_frame_transed_reg[8]_i_1_n_7 ;
  wire \control_frame_transed_reg[8]_i_1_n_8 ;
  wire \control_frame_transed_reg[8]_i_1_n_9 ;
  wire data_sel;
  wire data_sel_i_2_n_0;
  wire \fcs_error[0]_i_2_n_0 ;
  wire [63:0]fcs_error_reg;
  wire \fcs_error_reg[0]_i_1_n_0 ;
  wire \fcs_error_reg[0]_i_1_n_1 ;
  wire \fcs_error_reg[0]_i_1_n_10 ;
  wire \fcs_error_reg[0]_i_1_n_11 ;
  wire \fcs_error_reg[0]_i_1_n_12 ;
  wire \fcs_error_reg[0]_i_1_n_13 ;
  wire \fcs_error_reg[0]_i_1_n_14 ;
  wire \fcs_error_reg[0]_i_1_n_15 ;
  wire \fcs_error_reg[0]_i_1_n_2 ;
  wire \fcs_error_reg[0]_i_1_n_3 ;
  wire \fcs_error_reg[0]_i_1_n_4 ;
  wire \fcs_error_reg[0]_i_1_n_5 ;
  wire \fcs_error_reg[0]_i_1_n_6 ;
  wire \fcs_error_reg[0]_i_1_n_7 ;
  wire \fcs_error_reg[0]_i_1_n_8 ;
  wire \fcs_error_reg[0]_i_1_n_9 ;
  wire \fcs_error_reg[16]_i_1_n_0 ;
  wire \fcs_error_reg[16]_i_1_n_1 ;
  wire \fcs_error_reg[16]_i_1_n_10 ;
  wire \fcs_error_reg[16]_i_1_n_11 ;
  wire \fcs_error_reg[16]_i_1_n_12 ;
  wire \fcs_error_reg[16]_i_1_n_13 ;
  wire \fcs_error_reg[16]_i_1_n_14 ;
  wire \fcs_error_reg[16]_i_1_n_15 ;
  wire \fcs_error_reg[16]_i_1_n_2 ;
  wire \fcs_error_reg[16]_i_1_n_3 ;
  wire \fcs_error_reg[16]_i_1_n_4 ;
  wire \fcs_error_reg[16]_i_1_n_5 ;
  wire \fcs_error_reg[16]_i_1_n_6 ;
  wire \fcs_error_reg[16]_i_1_n_7 ;
  wire \fcs_error_reg[16]_i_1_n_8 ;
  wire \fcs_error_reg[16]_i_1_n_9 ;
  wire \fcs_error_reg[24]_i_1_n_0 ;
  wire \fcs_error_reg[24]_i_1_n_1 ;
  wire \fcs_error_reg[24]_i_1_n_10 ;
  wire \fcs_error_reg[24]_i_1_n_11 ;
  wire \fcs_error_reg[24]_i_1_n_12 ;
  wire \fcs_error_reg[24]_i_1_n_13 ;
  wire \fcs_error_reg[24]_i_1_n_14 ;
  wire \fcs_error_reg[24]_i_1_n_15 ;
  wire \fcs_error_reg[24]_i_1_n_2 ;
  wire \fcs_error_reg[24]_i_1_n_3 ;
  wire \fcs_error_reg[24]_i_1_n_4 ;
  wire \fcs_error_reg[24]_i_1_n_5 ;
  wire \fcs_error_reg[24]_i_1_n_6 ;
  wire \fcs_error_reg[24]_i_1_n_7 ;
  wire \fcs_error_reg[24]_i_1_n_8 ;
  wire \fcs_error_reg[24]_i_1_n_9 ;
  wire \fcs_error_reg[32]_i_1_n_0 ;
  wire \fcs_error_reg[32]_i_1_n_1 ;
  wire \fcs_error_reg[32]_i_1_n_10 ;
  wire \fcs_error_reg[32]_i_1_n_11 ;
  wire \fcs_error_reg[32]_i_1_n_12 ;
  wire \fcs_error_reg[32]_i_1_n_13 ;
  wire \fcs_error_reg[32]_i_1_n_14 ;
  wire \fcs_error_reg[32]_i_1_n_15 ;
  wire \fcs_error_reg[32]_i_1_n_2 ;
  wire \fcs_error_reg[32]_i_1_n_3 ;
  wire \fcs_error_reg[32]_i_1_n_4 ;
  wire \fcs_error_reg[32]_i_1_n_5 ;
  wire \fcs_error_reg[32]_i_1_n_6 ;
  wire \fcs_error_reg[32]_i_1_n_7 ;
  wire \fcs_error_reg[32]_i_1_n_8 ;
  wire \fcs_error_reg[32]_i_1_n_9 ;
  wire \fcs_error_reg[40]_i_1_n_0 ;
  wire \fcs_error_reg[40]_i_1_n_1 ;
  wire \fcs_error_reg[40]_i_1_n_10 ;
  wire \fcs_error_reg[40]_i_1_n_11 ;
  wire \fcs_error_reg[40]_i_1_n_12 ;
  wire \fcs_error_reg[40]_i_1_n_13 ;
  wire \fcs_error_reg[40]_i_1_n_14 ;
  wire \fcs_error_reg[40]_i_1_n_15 ;
  wire \fcs_error_reg[40]_i_1_n_2 ;
  wire \fcs_error_reg[40]_i_1_n_3 ;
  wire \fcs_error_reg[40]_i_1_n_4 ;
  wire \fcs_error_reg[40]_i_1_n_5 ;
  wire \fcs_error_reg[40]_i_1_n_6 ;
  wire \fcs_error_reg[40]_i_1_n_7 ;
  wire \fcs_error_reg[40]_i_1_n_8 ;
  wire \fcs_error_reg[40]_i_1_n_9 ;
  wire \fcs_error_reg[48]_i_1_n_0 ;
  wire \fcs_error_reg[48]_i_1_n_1 ;
  wire \fcs_error_reg[48]_i_1_n_10 ;
  wire \fcs_error_reg[48]_i_1_n_11 ;
  wire \fcs_error_reg[48]_i_1_n_12 ;
  wire \fcs_error_reg[48]_i_1_n_13 ;
  wire \fcs_error_reg[48]_i_1_n_14 ;
  wire \fcs_error_reg[48]_i_1_n_15 ;
  wire \fcs_error_reg[48]_i_1_n_2 ;
  wire \fcs_error_reg[48]_i_1_n_3 ;
  wire \fcs_error_reg[48]_i_1_n_4 ;
  wire \fcs_error_reg[48]_i_1_n_5 ;
  wire \fcs_error_reg[48]_i_1_n_6 ;
  wire \fcs_error_reg[48]_i_1_n_7 ;
  wire \fcs_error_reg[48]_i_1_n_8 ;
  wire \fcs_error_reg[48]_i_1_n_9 ;
  wire \fcs_error_reg[56]_i_1_n_1 ;
  wire \fcs_error_reg[56]_i_1_n_10 ;
  wire \fcs_error_reg[56]_i_1_n_11 ;
  wire \fcs_error_reg[56]_i_1_n_12 ;
  wire \fcs_error_reg[56]_i_1_n_13 ;
  wire \fcs_error_reg[56]_i_1_n_14 ;
  wire \fcs_error_reg[56]_i_1_n_15 ;
  wire \fcs_error_reg[56]_i_1_n_2 ;
  wire \fcs_error_reg[56]_i_1_n_3 ;
  wire \fcs_error_reg[56]_i_1_n_4 ;
  wire \fcs_error_reg[56]_i_1_n_5 ;
  wire \fcs_error_reg[56]_i_1_n_6 ;
  wire \fcs_error_reg[56]_i_1_n_7 ;
  wire \fcs_error_reg[56]_i_1_n_8 ;
  wire \fcs_error_reg[56]_i_1_n_9 ;
  wire \fcs_error_reg[8]_i_1_n_0 ;
  wire \fcs_error_reg[8]_i_1_n_1 ;
  wire \fcs_error_reg[8]_i_1_n_10 ;
  wire \fcs_error_reg[8]_i_1_n_11 ;
  wire \fcs_error_reg[8]_i_1_n_12 ;
  wire \fcs_error_reg[8]_i_1_n_13 ;
  wire \fcs_error_reg[8]_i_1_n_14 ;
  wire \fcs_error_reg[8]_i_1_n_15 ;
  wire \fcs_error_reg[8]_i_1_n_2 ;
  wire \fcs_error_reg[8]_i_1_n_3 ;
  wire \fcs_error_reg[8]_i_1_n_4 ;
  wire \fcs_error_reg[8]_i_1_n_5 ;
  wire \fcs_error_reg[8]_i_1_n_6 ;
  wire \fcs_error_reg[8]_i_1_n_7 ;
  wire \fcs_error_reg[8]_i_1_n_8 ;
  wire \fcs_error_reg[8]_i_1_n_9 ;
  wire \flow_control_config[31]_i_1_n_0 ;
  wire \flow_control_config[31]_i_2_n_0 ;
  wire \flow_control_config_reg_n_0_[0] ;
  wire \flow_control_config_reg_n_0_[10] ;
  wire \flow_control_config_reg_n_0_[11] ;
  wire \flow_control_config_reg_n_0_[12] ;
  wire \flow_control_config_reg_n_0_[13] ;
  wire \flow_control_config_reg_n_0_[14] ;
  wire \flow_control_config_reg_n_0_[15] ;
  wire \flow_control_config_reg_n_0_[16] ;
  wire \flow_control_config_reg_n_0_[17] ;
  wire \flow_control_config_reg_n_0_[18] ;
  wire \flow_control_config_reg_n_0_[19] ;
  wire \flow_control_config_reg_n_0_[1] ;
  wire \flow_control_config_reg_n_0_[20] ;
  wire \flow_control_config_reg_n_0_[21] ;
  wire \flow_control_config_reg_n_0_[22] ;
  wire \flow_control_config_reg_n_0_[23] ;
  wire \flow_control_config_reg_n_0_[24] ;
  wire \flow_control_config_reg_n_0_[25] ;
  wire \flow_control_config_reg_n_0_[26] ;
  wire \flow_control_config_reg_n_0_[27] ;
  wire \flow_control_config_reg_n_0_[28] ;
  wire \flow_control_config_reg_n_0_[29] ;
  wire \flow_control_config_reg_n_0_[2] ;
  wire \flow_control_config_reg_n_0_[31] ;
  wire \flow_control_config_reg_n_0_[3] ;
  wire \flow_control_config_reg_n_0_[4] ;
  wire \flow_control_config_reg_n_0_[5] ;
  wire \flow_control_config_reg_n_0_[6] ;
  wire \flow_control_config_reg_n_0_[7] ;
  wire \flow_control_config_reg_n_0_[8] ;
  wire \flow_control_config_reg_n_0_[9] ;
  wire \fragment_frame[0]_i_2_n_0 ;
  wire [63:0]fragment_frame_reg;
  wire \fragment_frame_reg[0]_i_1_n_0 ;
  wire \fragment_frame_reg[0]_i_1_n_1 ;
  wire \fragment_frame_reg[0]_i_1_n_10 ;
  wire \fragment_frame_reg[0]_i_1_n_11 ;
  wire \fragment_frame_reg[0]_i_1_n_12 ;
  wire \fragment_frame_reg[0]_i_1_n_13 ;
  wire \fragment_frame_reg[0]_i_1_n_14 ;
  wire \fragment_frame_reg[0]_i_1_n_15 ;
  wire \fragment_frame_reg[0]_i_1_n_2 ;
  wire \fragment_frame_reg[0]_i_1_n_3 ;
  wire \fragment_frame_reg[0]_i_1_n_4 ;
  wire \fragment_frame_reg[0]_i_1_n_5 ;
  wire \fragment_frame_reg[0]_i_1_n_6 ;
  wire \fragment_frame_reg[0]_i_1_n_7 ;
  wire \fragment_frame_reg[0]_i_1_n_8 ;
  wire \fragment_frame_reg[0]_i_1_n_9 ;
  wire \fragment_frame_reg[16]_i_1_n_0 ;
  wire \fragment_frame_reg[16]_i_1_n_1 ;
  wire \fragment_frame_reg[16]_i_1_n_10 ;
  wire \fragment_frame_reg[16]_i_1_n_11 ;
  wire \fragment_frame_reg[16]_i_1_n_12 ;
  wire \fragment_frame_reg[16]_i_1_n_13 ;
  wire \fragment_frame_reg[16]_i_1_n_14 ;
  wire \fragment_frame_reg[16]_i_1_n_15 ;
  wire \fragment_frame_reg[16]_i_1_n_2 ;
  wire \fragment_frame_reg[16]_i_1_n_3 ;
  wire \fragment_frame_reg[16]_i_1_n_4 ;
  wire \fragment_frame_reg[16]_i_1_n_5 ;
  wire \fragment_frame_reg[16]_i_1_n_6 ;
  wire \fragment_frame_reg[16]_i_1_n_7 ;
  wire \fragment_frame_reg[16]_i_1_n_8 ;
  wire \fragment_frame_reg[16]_i_1_n_9 ;
  wire \fragment_frame_reg[24]_i_1_n_0 ;
  wire \fragment_frame_reg[24]_i_1_n_1 ;
  wire \fragment_frame_reg[24]_i_1_n_10 ;
  wire \fragment_frame_reg[24]_i_1_n_11 ;
  wire \fragment_frame_reg[24]_i_1_n_12 ;
  wire \fragment_frame_reg[24]_i_1_n_13 ;
  wire \fragment_frame_reg[24]_i_1_n_14 ;
  wire \fragment_frame_reg[24]_i_1_n_15 ;
  wire \fragment_frame_reg[24]_i_1_n_2 ;
  wire \fragment_frame_reg[24]_i_1_n_3 ;
  wire \fragment_frame_reg[24]_i_1_n_4 ;
  wire \fragment_frame_reg[24]_i_1_n_5 ;
  wire \fragment_frame_reg[24]_i_1_n_6 ;
  wire \fragment_frame_reg[24]_i_1_n_7 ;
  wire \fragment_frame_reg[24]_i_1_n_8 ;
  wire \fragment_frame_reg[24]_i_1_n_9 ;
  wire \fragment_frame_reg[32]_i_1_n_0 ;
  wire \fragment_frame_reg[32]_i_1_n_1 ;
  wire \fragment_frame_reg[32]_i_1_n_10 ;
  wire \fragment_frame_reg[32]_i_1_n_11 ;
  wire \fragment_frame_reg[32]_i_1_n_12 ;
  wire \fragment_frame_reg[32]_i_1_n_13 ;
  wire \fragment_frame_reg[32]_i_1_n_14 ;
  wire \fragment_frame_reg[32]_i_1_n_15 ;
  wire \fragment_frame_reg[32]_i_1_n_2 ;
  wire \fragment_frame_reg[32]_i_1_n_3 ;
  wire \fragment_frame_reg[32]_i_1_n_4 ;
  wire \fragment_frame_reg[32]_i_1_n_5 ;
  wire \fragment_frame_reg[32]_i_1_n_6 ;
  wire \fragment_frame_reg[32]_i_1_n_7 ;
  wire \fragment_frame_reg[32]_i_1_n_8 ;
  wire \fragment_frame_reg[32]_i_1_n_9 ;
  wire \fragment_frame_reg[40]_i_1_n_0 ;
  wire \fragment_frame_reg[40]_i_1_n_1 ;
  wire \fragment_frame_reg[40]_i_1_n_10 ;
  wire \fragment_frame_reg[40]_i_1_n_11 ;
  wire \fragment_frame_reg[40]_i_1_n_12 ;
  wire \fragment_frame_reg[40]_i_1_n_13 ;
  wire \fragment_frame_reg[40]_i_1_n_14 ;
  wire \fragment_frame_reg[40]_i_1_n_15 ;
  wire \fragment_frame_reg[40]_i_1_n_2 ;
  wire \fragment_frame_reg[40]_i_1_n_3 ;
  wire \fragment_frame_reg[40]_i_1_n_4 ;
  wire \fragment_frame_reg[40]_i_1_n_5 ;
  wire \fragment_frame_reg[40]_i_1_n_6 ;
  wire \fragment_frame_reg[40]_i_1_n_7 ;
  wire \fragment_frame_reg[40]_i_1_n_8 ;
  wire \fragment_frame_reg[40]_i_1_n_9 ;
  wire \fragment_frame_reg[48]_i_1_n_0 ;
  wire \fragment_frame_reg[48]_i_1_n_1 ;
  wire \fragment_frame_reg[48]_i_1_n_10 ;
  wire \fragment_frame_reg[48]_i_1_n_11 ;
  wire \fragment_frame_reg[48]_i_1_n_12 ;
  wire \fragment_frame_reg[48]_i_1_n_13 ;
  wire \fragment_frame_reg[48]_i_1_n_14 ;
  wire \fragment_frame_reg[48]_i_1_n_15 ;
  wire \fragment_frame_reg[48]_i_1_n_2 ;
  wire \fragment_frame_reg[48]_i_1_n_3 ;
  wire \fragment_frame_reg[48]_i_1_n_4 ;
  wire \fragment_frame_reg[48]_i_1_n_5 ;
  wire \fragment_frame_reg[48]_i_1_n_6 ;
  wire \fragment_frame_reg[48]_i_1_n_7 ;
  wire \fragment_frame_reg[48]_i_1_n_8 ;
  wire \fragment_frame_reg[48]_i_1_n_9 ;
  wire \fragment_frame_reg[56]_i_1_n_1 ;
  wire \fragment_frame_reg[56]_i_1_n_10 ;
  wire \fragment_frame_reg[56]_i_1_n_11 ;
  wire \fragment_frame_reg[56]_i_1_n_12 ;
  wire \fragment_frame_reg[56]_i_1_n_13 ;
  wire \fragment_frame_reg[56]_i_1_n_14 ;
  wire \fragment_frame_reg[56]_i_1_n_15 ;
  wire \fragment_frame_reg[56]_i_1_n_2 ;
  wire \fragment_frame_reg[56]_i_1_n_3 ;
  wire \fragment_frame_reg[56]_i_1_n_4 ;
  wire \fragment_frame_reg[56]_i_1_n_5 ;
  wire \fragment_frame_reg[56]_i_1_n_6 ;
  wire \fragment_frame_reg[56]_i_1_n_7 ;
  wire \fragment_frame_reg[56]_i_1_n_8 ;
  wire \fragment_frame_reg[56]_i_1_n_9 ;
  wire \fragment_frame_reg[8]_i_1_n_0 ;
  wire \fragment_frame_reg[8]_i_1_n_1 ;
  wire \fragment_frame_reg[8]_i_1_n_10 ;
  wire \fragment_frame_reg[8]_i_1_n_11 ;
  wire \fragment_frame_reg[8]_i_1_n_12 ;
  wire \fragment_frame_reg[8]_i_1_n_13 ;
  wire \fragment_frame_reg[8]_i_1_n_14 ;
  wire \fragment_frame_reg[8]_i_1_n_15 ;
  wire \fragment_frame_reg[8]_i_1_n_2 ;
  wire \fragment_frame_reg[8]_i_1_n_3 ;
  wire \fragment_frame_reg[8]_i_1_n_4 ;
  wire \fragment_frame_reg[8]_i_1_n_5 ;
  wire \fragment_frame_reg[8]_i_1_n_6 ;
  wire \fragment_frame_reg[8]_i_1_n_7 ;
  wire \fragment_frame_reg[8]_i_1_n_8 ;
  wire \fragment_frame_reg[8]_i_1_n_9 ;
  wire \frame_1024_max_good[0]_i_2_n_0 ;
  wire [63:0]frame_1024_max_good_reg;
  wire \frame_1024_max_good_reg[0]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[0]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[16]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[24]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[32]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[40]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[48]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[56]_i_1_n_9 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_0 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_1 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_10 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_11 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_12 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_13 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_14 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_15 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_2 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_3 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_4 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_5 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_6 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_7 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_8 ;
  wire \frame_1024_max_good_reg[8]_i_1_n_9 ;
  wire \frame_1024_max_transed[0]_i_2_n_0 ;
  wire [63:0]frame_1024_max_transed_reg;
  wire \frame_1024_max_transed_reg[0]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[0]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[16]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[24]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[32]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[40]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[48]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[56]_i_1_n_9 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_0 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_1 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_10 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_11 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_12 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_13 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_14 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_15 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_2 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_3 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_4 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_5 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_6 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_7 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_8 ;
  wire \frame_1024_max_transed_reg[8]_i_1_n_9 ;
  wire \frame_128_255_good[0]_i_2_n_0 ;
  wire [63:0]frame_128_255_good_reg;
  wire \frame_128_255_good_reg[0]_i_1_n_0 ;
  wire \frame_128_255_good_reg[0]_i_1_n_1 ;
  wire \frame_128_255_good_reg[0]_i_1_n_10 ;
  wire \frame_128_255_good_reg[0]_i_1_n_11 ;
  wire \frame_128_255_good_reg[0]_i_1_n_12 ;
  wire \frame_128_255_good_reg[0]_i_1_n_13 ;
  wire \frame_128_255_good_reg[0]_i_1_n_14 ;
  wire \frame_128_255_good_reg[0]_i_1_n_15 ;
  wire \frame_128_255_good_reg[0]_i_1_n_2 ;
  wire \frame_128_255_good_reg[0]_i_1_n_3 ;
  wire \frame_128_255_good_reg[0]_i_1_n_4 ;
  wire \frame_128_255_good_reg[0]_i_1_n_5 ;
  wire \frame_128_255_good_reg[0]_i_1_n_6 ;
  wire \frame_128_255_good_reg[0]_i_1_n_7 ;
  wire \frame_128_255_good_reg[0]_i_1_n_8 ;
  wire \frame_128_255_good_reg[0]_i_1_n_9 ;
  wire \frame_128_255_good_reg[16]_i_1_n_0 ;
  wire \frame_128_255_good_reg[16]_i_1_n_1 ;
  wire \frame_128_255_good_reg[16]_i_1_n_10 ;
  wire \frame_128_255_good_reg[16]_i_1_n_11 ;
  wire \frame_128_255_good_reg[16]_i_1_n_12 ;
  wire \frame_128_255_good_reg[16]_i_1_n_13 ;
  wire \frame_128_255_good_reg[16]_i_1_n_14 ;
  wire \frame_128_255_good_reg[16]_i_1_n_15 ;
  wire \frame_128_255_good_reg[16]_i_1_n_2 ;
  wire \frame_128_255_good_reg[16]_i_1_n_3 ;
  wire \frame_128_255_good_reg[16]_i_1_n_4 ;
  wire \frame_128_255_good_reg[16]_i_1_n_5 ;
  wire \frame_128_255_good_reg[16]_i_1_n_6 ;
  wire \frame_128_255_good_reg[16]_i_1_n_7 ;
  wire \frame_128_255_good_reg[16]_i_1_n_8 ;
  wire \frame_128_255_good_reg[16]_i_1_n_9 ;
  wire \frame_128_255_good_reg[24]_i_1_n_0 ;
  wire \frame_128_255_good_reg[24]_i_1_n_1 ;
  wire \frame_128_255_good_reg[24]_i_1_n_10 ;
  wire \frame_128_255_good_reg[24]_i_1_n_11 ;
  wire \frame_128_255_good_reg[24]_i_1_n_12 ;
  wire \frame_128_255_good_reg[24]_i_1_n_13 ;
  wire \frame_128_255_good_reg[24]_i_1_n_14 ;
  wire \frame_128_255_good_reg[24]_i_1_n_15 ;
  wire \frame_128_255_good_reg[24]_i_1_n_2 ;
  wire \frame_128_255_good_reg[24]_i_1_n_3 ;
  wire \frame_128_255_good_reg[24]_i_1_n_4 ;
  wire \frame_128_255_good_reg[24]_i_1_n_5 ;
  wire \frame_128_255_good_reg[24]_i_1_n_6 ;
  wire \frame_128_255_good_reg[24]_i_1_n_7 ;
  wire \frame_128_255_good_reg[24]_i_1_n_8 ;
  wire \frame_128_255_good_reg[24]_i_1_n_9 ;
  wire \frame_128_255_good_reg[32]_i_1_n_0 ;
  wire \frame_128_255_good_reg[32]_i_1_n_1 ;
  wire \frame_128_255_good_reg[32]_i_1_n_10 ;
  wire \frame_128_255_good_reg[32]_i_1_n_11 ;
  wire \frame_128_255_good_reg[32]_i_1_n_12 ;
  wire \frame_128_255_good_reg[32]_i_1_n_13 ;
  wire \frame_128_255_good_reg[32]_i_1_n_14 ;
  wire \frame_128_255_good_reg[32]_i_1_n_15 ;
  wire \frame_128_255_good_reg[32]_i_1_n_2 ;
  wire \frame_128_255_good_reg[32]_i_1_n_3 ;
  wire \frame_128_255_good_reg[32]_i_1_n_4 ;
  wire \frame_128_255_good_reg[32]_i_1_n_5 ;
  wire \frame_128_255_good_reg[32]_i_1_n_6 ;
  wire \frame_128_255_good_reg[32]_i_1_n_7 ;
  wire \frame_128_255_good_reg[32]_i_1_n_8 ;
  wire \frame_128_255_good_reg[32]_i_1_n_9 ;
  wire \frame_128_255_good_reg[40]_i_1_n_0 ;
  wire \frame_128_255_good_reg[40]_i_1_n_1 ;
  wire \frame_128_255_good_reg[40]_i_1_n_10 ;
  wire \frame_128_255_good_reg[40]_i_1_n_11 ;
  wire \frame_128_255_good_reg[40]_i_1_n_12 ;
  wire \frame_128_255_good_reg[40]_i_1_n_13 ;
  wire \frame_128_255_good_reg[40]_i_1_n_14 ;
  wire \frame_128_255_good_reg[40]_i_1_n_15 ;
  wire \frame_128_255_good_reg[40]_i_1_n_2 ;
  wire \frame_128_255_good_reg[40]_i_1_n_3 ;
  wire \frame_128_255_good_reg[40]_i_1_n_4 ;
  wire \frame_128_255_good_reg[40]_i_1_n_5 ;
  wire \frame_128_255_good_reg[40]_i_1_n_6 ;
  wire \frame_128_255_good_reg[40]_i_1_n_7 ;
  wire \frame_128_255_good_reg[40]_i_1_n_8 ;
  wire \frame_128_255_good_reg[40]_i_1_n_9 ;
  wire \frame_128_255_good_reg[48]_i_1_n_0 ;
  wire \frame_128_255_good_reg[48]_i_1_n_1 ;
  wire \frame_128_255_good_reg[48]_i_1_n_10 ;
  wire \frame_128_255_good_reg[48]_i_1_n_11 ;
  wire \frame_128_255_good_reg[48]_i_1_n_12 ;
  wire \frame_128_255_good_reg[48]_i_1_n_13 ;
  wire \frame_128_255_good_reg[48]_i_1_n_14 ;
  wire \frame_128_255_good_reg[48]_i_1_n_15 ;
  wire \frame_128_255_good_reg[48]_i_1_n_2 ;
  wire \frame_128_255_good_reg[48]_i_1_n_3 ;
  wire \frame_128_255_good_reg[48]_i_1_n_4 ;
  wire \frame_128_255_good_reg[48]_i_1_n_5 ;
  wire \frame_128_255_good_reg[48]_i_1_n_6 ;
  wire \frame_128_255_good_reg[48]_i_1_n_7 ;
  wire \frame_128_255_good_reg[48]_i_1_n_8 ;
  wire \frame_128_255_good_reg[48]_i_1_n_9 ;
  wire \frame_128_255_good_reg[56]_i_1_n_1 ;
  wire \frame_128_255_good_reg[56]_i_1_n_10 ;
  wire \frame_128_255_good_reg[56]_i_1_n_11 ;
  wire \frame_128_255_good_reg[56]_i_1_n_12 ;
  wire \frame_128_255_good_reg[56]_i_1_n_13 ;
  wire \frame_128_255_good_reg[56]_i_1_n_14 ;
  wire \frame_128_255_good_reg[56]_i_1_n_15 ;
  wire \frame_128_255_good_reg[56]_i_1_n_2 ;
  wire \frame_128_255_good_reg[56]_i_1_n_3 ;
  wire \frame_128_255_good_reg[56]_i_1_n_4 ;
  wire \frame_128_255_good_reg[56]_i_1_n_5 ;
  wire \frame_128_255_good_reg[56]_i_1_n_6 ;
  wire \frame_128_255_good_reg[56]_i_1_n_7 ;
  wire \frame_128_255_good_reg[56]_i_1_n_8 ;
  wire \frame_128_255_good_reg[56]_i_1_n_9 ;
  wire \frame_128_255_good_reg[8]_i_1_n_0 ;
  wire \frame_128_255_good_reg[8]_i_1_n_1 ;
  wire \frame_128_255_good_reg[8]_i_1_n_10 ;
  wire \frame_128_255_good_reg[8]_i_1_n_11 ;
  wire \frame_128_255_good_reg[8]_i_1_n_12 ;
  wire \frame_128_255_good_reg[8]_i_1_n_13 ;
  wire \frame_128_255_good_reg[8]_i_1_n_14 ;
  wire \frame_128_255_good_reg[8]_i_1_n_15 ;
  wire \frame_128_255_good_reg[8]_i_1_n_2 ;
  wire \frame_128_255_good_reg[8]_i_1_n_3 ;
  wire \frame_128_255_good_reg[8]_i_1_n_4 ;
  wire \frame_128_255_good_reg[8]_i_1_n_5 ;
  wire \frame_128_255_good_reg[8]_i_1_n_6 ;
  wire \frame_128_255_good_reg[8]_i_1_n_7 ;
  wire \frame_128_255_good_reg[8]_i_1_n_8 ;
  wire \frame_128_255_good_reg[8]_i_1_n_9 ;
  wire \frame_128_255_transed[0]_i_2_n_0 ;
  wire [63:0]frame_128_255_transed_reg;
  wire \frame_128_255_transed_reg[0]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[0]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[16]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[24]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[32]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[40]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[48]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[56]_i_1_n_9 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_0 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_1 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_10 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_11 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_12 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_13 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_14 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_15 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_2 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_3 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_4 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_5 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_6 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_7 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_8 ;
  wire \frame_128_255_transed_reg[8]_i_1_n_9 ;
  wire \frame_256_511_good[0]_i_2_n_0 ;
  wire [63:0]frame_256_511_good_reg;
  wire \frame_256_511_good_reg[0]_i_1_n_0 ;
  wire \frame_256_511_good_reg[0]_i_1_n_1 ;
  wire \frame_256_511_good_reg[0]_i_1_n_10 ;
  wire \frame_256_511_good_reg[0]_i_1_n_11 ;
  wire \frame_256_511_good_reg[0]_i_1_n_12 ;
  wire \frame_256_511_good_reg[0]_i_1_n_13 ;
  wire \frame_256_511_good_reg[0]_i_1_n_14 ;
  wire \frame_256_511_good_reg[0]_i_1_n_15 ;
  wire \frame_256_511_good_reg[0]_i_1_n_2 ;
  wire \frame_256_511_good_reg[0]_i_1_n_3 ;
  wire \frame_256_511_good_reg[0]_i_1_n_4 ;
  wire \frame_256_511_good_reg[0]_i_1_n_5 ;
  wire \frame_256_511_good_reg[0]_i_1_n_6 ;
  wire \frame_256_511_good_reg[0]_i_1_n_7 ;
  wire \frame_256_511_good_reg[0]_i_1_n_8 ;
  wire \frame_256_511_good_reg[0]_i_1_n_9 ;
  wire \frame_256_511_good_reg[16]_i_1_n_0 ;
  wire \frame_256_511_good_reg[16]_i_1_n_1 ;
  wire \frame_256_511_good_reg[16]_i_1_n_10 ;
  wire \frame_256_511_good_reg[16]_i_1_n_11 ;
  wire \frame_256_511_good_reg[16]_i_1_n_12 ;
  wire \frame_256_511_good_reg[16]_i_1_n_13 ;
  wire \frame_256_511_good_reg[16]_i_1_n_14 ;
  wire \frame_256_511_good_reg[16]_i_1_n_15 ;
  wire \frame_256_511_good_reg[16]_i_1_n_2 ;
  wire \frame_256_511_good_reg[16]_i_1_n_3 ;
  wire \frame_256_511_good_reg[16]_i_1_n_4 ;
  wire \frame_256_511_good_reg[16]_i_1_n_5 ;
  wire \frame_256_511_good_reg[16]_i_1_n_6 ;
  wire \frame_256_511_good_reg[16]_i_1_n_7 ;
  wire \frame_256_511_good_reg[16]_i_1_n_8 ;
  wire \frame_256_511_good_reg[16]_i_1_n_9 ;
  wire \frame_256_511_good_reg[24]_i_1_n_0 ;
  wire \frame_256_511_good_reg[24]_i_1_n_1 ;
  wire \frame_256_511_good_reg[24]_i_1_n_10 ;
  wire \frame_256_511_good_reg[24]_i_1_n_11 ;
  wire \frame_256_511_good_reg[24]_i_1_n_12 ;
  wire \frame_256_511_good_reg[24]_i_1_n_13 ;
  wire \frame_256_511_good_reg[24]_i_1_n_14 ;
  wire \frame_256_511_good_reg[24]_i_1_n_15 ;
  wire \frame_256_511_good_reg[24]_i_1_n_2 ;
  wire \frame_256_511_good_reg[24]_i_1_n_3 ;
  wire \frame_256_511_good_reg[24]_i_1_n_4 ;
  wire \frame_256_511_good_reg[24]_i_1_n_5 ;
  wire \frame_256_511_good_reg[24]_i_1_n_6 ;
  wire \frame_256_511_good_reg[24]_i_1_n_7 ;
  wire \frame_256_511_good_reg[24]_i_1_n_8 ;
  wire \frame_256_511_good_reg[24]_i_1_n_9 ;
  wire \frame_256_511_good_reg[32]_i_1_n_0 ;
  wire \frame_256_511_good_reg[32]_i_1_n_1 ;
  wire \frame_256_511_good_reg[32]_i_1_n_10 ;
  wire \frame_256_511_good_reg[32]_i_1_n_11 ;
  wire \frame_256_511_good_reg[32]_i_1_n_12 ;
  wire \frame_256_511_good_reg[32]_i_1_n_13 ;
  wire \frame_256_511_good_reg[32]_i_1_n_14 ;
  wire \frame_256_511_good_reg[32]_i_1_n_15 ;
  wire \frame_256_511_good_reg[32]_i_1_n_2 ;
  wire \frame_256_511_good_reg[32]_i_1_n_3 ;
  wire \frame_256_511_good_reg[32]_i_1_n_4 ;
  wire \frame_256_511_good_reg[32]_i_1_n_5 ;
  wire \frame_256_511_good_reg[32]_i_1_n_6 ;
  wire \frame_256_511_good_reg[32]_i_1_n_7 ;
  wire \frame_256_511_good_reg[32]_i_1_n_8 ;
  wire \frame_256_511_good_reg[32]_i_1_n_9 ;
  wire \frame_256_511_good_reg[40]_i_1_n_0 ;
  wire \frame_256_511_good_reg[40]_i_1_n_1 ;
  wire \frame_256_511_good_reg[40]_i_1_n_10 ;
  wire \frame_256_511_good_reg[40]_i_1_n_11 ;
  wire \frame_256_511_good_reg[40]_i_1_n_12 ;
  wire \frame_256_511_good_reg[40]_i_1_n_13 ;
  wire \frame_256_511_good_reg[40]_i_1_n_14 ;
  wire \frame_256_511_good_reg[40]_i_1_n_15 ;
  wire \frame_256_511_good_reg[40]_i_1_n_2 ;
  wire \frame_256_511_good_reg[40]_i_1_n_3 ;
  wire \frame_256_511_good_reg[40]_i_1_n_4 ;
  wire \frame_256_511_good_reg[40]_i_1_n_5 ;
  wire \frame_256_511_good_reg[40]_i_1_n_6 ;
  wire \frame_256_511_good_reg[40]_i_1_n_7 ;
  wire \frame_256_511_good_reg[40]_i_1_n_8 ;
  wire \frame_256_511_good_reg[40]_i_1_n_9 ;
  wire \frame_256_511_good_reg[48]_i_1_n_0 ;
  wire \frame_256_511_good_reg[48]_i_1_n_1 ;
  wire \frame_256_511_good_reg[48]_i_1_n_10 ;
  wire \frame_256_511_good_reg[48]_i_1_n_11 ;
  wire \frame_256_511_good_reg[48]_i_1_n_12 ;
  wire \frame_256_511_good_reg[48]_i_1_n_13 ;
  wire \frame_256_511_good_reg[48]_i_1_n_14 ;
  wire \frame_256_511_good_reg[48]_i_1_n_15 ;
  wire \frame_256_511_good_reg[48]_i_1_n_2 ;
  wire \frame_256_511_good_reg[48]_i_1_n_3 ;
  wire \frame_256_511_good_reg[48]_i_1_n_4 ;
  wire \frame_256_511_good_reg[48]_i_1_n_5 ;
  wire \frame_256_511_good_reg[48]_i_1_n_6 ;
  wire \frame_256_511_good_reg[48]_i_1_n_7 ;
  wire \frame_256_511_good_reg[48]_i_1_n_8 ;
  wire \frame_256_511_good_reg[48]_i_1_n_9 ;
  wire \frame_256_511_good_reg[56]_i_1_n_1 ;
  wire \frame_256_511_good_reg[56]_i_1_n_10 ;
  wire \frame_256_511_good_reg[56]_i_1_n_11 ;
  wire \frame_256_511_good_reg[56]_i_1_n_12 ;
  wire \frame_256_511_good_reg[56]_i_1_n_13 ;
  wire \frame_256_511_good_reg[56]_i_1_n_14 ;
  wire \frame_256_511_good_reg[56]_i_1_n_15 ;
  wire \frame_256_511_good_reg[56]_i_1_n_2 ;
  wire \frame_256_511_good_reg[56]_i_1_n_3 ;
  wire \frame_256_511_good_reg[56]_i_1_n_4 ;
  wire \frame_256_511_good_reg[56]_i_1_n_5 ;
  wire \frame_256_511_good_reg[56]_i_1_n_6 ;
  wire \frame_256_511_good_reg[56]_i_1_n_7 ;
  wire \frame_256_511_good_reg[56]_i_1_n_8 ;
  wire \frame_256_511_good_reg[56]_i_1_n_9 ;
  wire \frame_256_511_good_reg[8]_i_1_n_0 ;
  wire \frame_256_511_good_reg[8]_i_1_n_1 ;
  wire \frame_256_511_good_reg[8]_i_1_n_10 ;
  wire \frame_256_511_good_reg[8]_i_1_n_11 ;
  wire \frame_256_511_good_reg[8]_i_1_n_12 ;
  wire \frame_256_511_good_reg[8]_i_1_n_13 ;
  wire \frame_256_511_good_reg[8]_i_1_n_14 ;
  wire \frame_256_511_good_reg[8]_i_1_n_15 ;
  wire \frame_256_511_good_reg[8]_i_1_n_2 ;
  wire \frame_256_511_good_reg[8]_i_1_n_3 ;
  wire \frame_256_511_good_reg[8]_i_1_n_4 ;
  wire \frame_256_511_good_reg[8]_i_1_n_5 ;
  wire \frame_256_511_good_reg[8]_i_1_n_6 ;
  wire \frame_256_511_good_reg[8]_i_1_n_7 ;
  wire \frame_256_511_good_reg[8]_i_1_n_8 ;
  wire \frame_256_511_good_reg[8]_i_1_n_9 ;
  wire \frame_256_511_transed[0]_i_2_n_0 ;
  wire [63:0]frame_256_511_transed_reg;
  wire \frame_256_511_transed_reg[0]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[0]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[16]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[24]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[32]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[40]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[48]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[56]_i_1_n_9 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_0 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_1 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_10 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_11 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_12 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_13 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_14 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_15 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_2 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_3 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_4 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_5 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_6 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_7 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_8 ;
  wire \frame_256_511_transed_reg[8]_i_1_n_9 ;
  wire \frame_512_1023_good[0]_i_2_n_0 ;
  wire [63:0]frame_512_1023_good_reg;
  wire \frame_512_1023_good_reg[0]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[0]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[16]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[24]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[32]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[40]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[48]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[56]_i_1_n_9 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_0 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_1 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_10 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_11 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_12 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_13 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_14 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_15 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_2 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_3 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_4 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_5 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_6 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_7 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_8 ;
  wire \frame_512_1023_good_reg[8]_i_1_n_9 ;
  wire \frame_512_1023_transed[0]_i_2_n_0 ;
  wire [63:0]frame_512_1023_transed_reg;
  wire \frame_512_1023_transed_reg[0]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[0]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[16]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[24]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[32]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[40]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[48]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[56]_i_1_n_9 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_0 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_1 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_10 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_11 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_12 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_13 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_14 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_15 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_2 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_3 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_4 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_5 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_6 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_7 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_8 ;
  wire \frame_512_1023_transed_reg[8]_i_1_n_9 ;
  wire \frame_64_good[0]_i_2_n_0 ;
  wire [63:0]frame_64_good_reg;
  wire \frame_64_good_reg[0]_i_1_n_0 ;
  wire \frame_64_good_reg[0]_i_1_n_1 ;
  wire \frame_64_good_reg[0]_i_1_n_10 ;
  wire \frame_64_good_reg[0]_i_1_n_11 ;
  wire \frame_64_good_reg[0]_i_1_n_12 ;
  wire \frame_64_good_reg[0]_i_1_n_13 ;
  wire \frame_64_good_reg[0]_i_1_n_14 ;
  wire \frame_64_good_reg[0]_i_1_n_15 ;
  wire \frame_64_good_reg[0]_i_1_n_2 ;
  wire \frame_64_good_reg[0]_i_1_n_3 ;
  wire \frame_64_good_reg[0]_i_1_n_4 ;
  wire \frame_64_good_reg[0]_i_1_n_5 ;
  wire \frame_64_good_reg[0]_i_1_n_6 ;
  wire \frame_64_good_reg[0]_i_1_n_7 ;
  wire \frame_64_good_reg[0]_i_1_n_8 ;
  wire \frame_64_good_reg[0]_i_1_n_9 ;
  wire \frame_64_good_reg[16]_i_1_n_0 ;
  wire \frame_64_good_reg[16]_i_1_n_1 ;
  wire \frame_64_good_reg[16]_i_1_n_10 ;
  wire \frame_64_good_reg[16]_i_1_n_11 ;
  wire \frame_64_good_reg[16]_i_1_n_12 ;
  wire \frame_64_good_reg[16]_i_1_n_13 ;
  wire \frame_64_good_reg[16]_i_1_n_14 ;
  wire \frame_64_good_reg[16]_i_1_n_15 ;
  wire \frame_64_good_reg[16]_i_1_n_2 ;
  wire \frame_64_good_reg[16]_i_1_n_3 ;
  wire \frame_64_good_reg[16]_i_1_n_4 ;
  wire \frame_64_good_reg[16]_i_1_n_5 ;
  wire \frame_64_good_reg[16]_i_1_n_6 ;
  wire \frame_64_good_reg[16]_i_1_n_7 ;
  wire \frame_64_good_reg[16]_i_1_n_8 ;
  wire \frame_64_good_reg[16]_i_1_n_9 ;
  wire \frame_64_good_reg[24]_i_1_n_0 ;
  wire \frame_64_good_reg[24]_i_1_n_1 ;
  wire \frame_64_good_reg[24]_i_1_n_10 ;
  wire \frame_64_good_reg[24]_i_1_n_11 ;
  wire \frame_64_good_reg[24]_i_1_n_12 ;
  wire \frame_64_good_reg[24]_i_1_n_13 ;
  wire \frame_64_good_reg[24]_i_1_n_14 ;
  wire \frame_64_good_reg[24]_i_1_n_15 ;
  wire \frame_64_good_reg[24]_i_1_n_2 ;
  wire \frame_64_good_reg[24]_i_1_n_3 ;
  wire \frame_64_good_reg[24]_i_1_n_4 ;
  wire \frame_64_good_reg[24]_i_1_n_5 ;
  wire \frame_64_good_reg[24]_i_1_n_6 ;
  wire \frame_64_good_reg[24]_i_1_n_7 ;
  wire \frame_64_good_reg[24]_i_1_n_8 ;
  wire \frame_64_good_reg[24]_i_1_n_9 ;
  wire \frame_64_good_reg[32]_i_1_n_0 ;
  wire \frame_64_good_reg[32]_i_1_n_1 ;
  wire \frame_64_good_reg[32]_i_1_n_10 ;
  wire \frame_64_good_reg[32]_i_1_n_11 ;
  wire \frame_64_good_reg[32]_i_1_n_12 ;
  wire \frame_64_good_reg[32]_i_1_n_13 ;
  wire \frame_64_good_reg[32]_i_1_n_14 ;
  wire \frame_64_good_reg[32]_i_1_n_15 ;
  wire \frame_64_good_reg[32]_i_1_n_2 ;
  wire \frame_64_good_reg[32]_i_1_n_3 ;
  wire \frame_64_good_reg[32]_i_1_n_4 ;
  wire \frame_64_good_reg[32]_i_1_n_5 ;
  wire \frame_64_good_reg[32]_i_1_n_6 ;
  wire \frame_64_good_reg[32]_i_1_n_7 ;
  wire \frame_64_good_reg[32]_i_1_n_8 ;
  wire \frame_64_good_reg[32]_i_1_n_9 ;
  wire \frame_64_good_reg[40]_i_1_n_0 ;
  wire \frame_64_good_reg[40]_i_1_n_1 ;
  wire \frame_64_good_reg[40]_i_1_n_10 ;
  wire \frame_64_good_reg[40]_i_1_n_11 ;
  wire \frame_64_good_reg[40]_i_1_n_12 ;
  wire \frame_64_good_reg[40]_i_1_n_13 ;
  wire \frame_64_good_reg[40]_i_1_n_14 ;
  wire \frame_64_good_reg[40]_i_1_n_15 ;
  wire \frame_64_good_reg[40]_i_1_n_2 ;
  wire \frame_64_good_reg[40]_i_1_n_3 ;
  wire \frame_64_good_reg[40]_i_1_n_4 ;
  wire \frame_64_good_reg[40]_i_1_n_5 ;
  wire \frame_64_good_reg[40]_i_1_n_6 ;
  wire \frame_64_good_reg[40]_i_1_n_7 ;
  wire \frame_64_good_reg[40]_i_1_n_8 ;
  wire \frame_64_good_reg[40]_i_1_n_9 ;
  wire \frame_64_good_reg[48]_i_1_n_0 ;
  wire \frame_64_good_reg[48]_i_1_n_1 ;
  wire \frame_64_good_reg[48]_i_1_n_10 ;
  wire \frame_64_good_reg[48]_i_1_n_11 ;
  wire \frame_64_good_reg[48]_i_1_n_12 ;
  wire \frame_64_good_reg[48]_i_1_n_13 ;
  wire \frame_64_good_reg[48]_i_1_n_14 ;
  wire \frame_64_good_reg[48]_i_1_n_15 ;
  wire \frame_64_good_reg[48]_i_1_n_2 ;
  wire \frame_64_good_reg[48]_i_1_n_3 ;
  wire \frame_64_good_reg[48]_i_1_n_4 ;
  wire \frame_64_good_reg[48]_i_1_n_5 ;
  wire \frame_64_good_reg[48]_i_1_n_6 ;
  wire \frame_64_good_reg[48]_i_1_n_7 ;
  wire \frame_64_good_reg[48]_i_1_n_8 ;
  wire \frame_64_good_reg[48]_i_1_n_9 ;
  wire \frame_64_good_reg[56]_i_1_n_1 ;
  wire \frame_64_good_reg[56]_i_1_n_10 ;
  wire \frame_64_good_reg[56]_i_1_n_11 ;
  wire \frame_64_good_reg[56]_i_1_n_12 ;
  wire \frame_64_good_reg[56]_i_1_n_13 ;
  wire \frame_64_good_reg[56]_i_1_n_14 ;
  wire \frame_64_good_reg[56]_i_1_n_15 ;
  wire \frame_64_good_reg[56]_i_1_n_2 ;
  wire \frame_64_good_reg[56]_i_1_n_3 ;
  wire \frame_64_good_reg[56]_i_1_n_4 ;
  wire \frame_64_good_reg[56]_i_1_n_5 ;
  wire \frame_64_good_reg[56]_i_1_n_6 ;
  wire \frame_64_good_reg[56]_i_1_n_7 ;
  wire \frame_64_good_reg[56]_i_1_n_8 ;
  wire \frame_64_good_reg[56]_i_1_n_9 ;
  wire \frame_64_good_reg[8]_i_1_n_0 ;
  wire \frame_64_good_reg[8]_i_1_n_1 ;
  wire \frame_64_good_reg[8]_i_1_n_10 ;
  wire \frame_64_good_reg[8]_i_1_n_11 ;
  wire \frame_64_good_reg[8]_i_1_n_12 ;
  wire \frame_64_good_reg[8]_i_1_n_13 ;
  wire \frame_64_good_reg[8]_i_1_n_14 ;
  wire \frame_64_good_reg[8]_i_1_n_15 ;
  wire \frame_64_good_reg[8]_i_1_n_2 ;
  wire \frame_64_good_reg[8]_i_1_n_3 ;
  wire \frame_64_good_reg[8]_i_1_n_4 ;
  wire \frame_64_good_reg[8]_i_1_n_5 ;
  wire \frame_64_good_reg[8]_i_1_n_6 ;
  wire \frame_64_good_reg[8]_i_1_n_7 ;
  wire \frame_64_good_reg[8]_i_1_n_8 ;
  wire \frame_64_good_reg[8]_i_1_n_9 ;
  wire \frame_64_transed[0]_i_2_n_0 ;
  wire [63:0]frame_64_transed_reg;
  wire \frame_64_transed_reg[0]_i_1_n_0 ;
  wire \frame_64_transed_reg[0]_i_1_n_1 ;
  wire \frame_64_transed_reg[0]_i_1_n_10 ;
  wire \frame_64_transed_reg[0]_i_1_n_11 ;
  wire \frame_64_transed_reg[0]_i_1_n_12 ;
  wire \frame_64_transed_reg[0]_i_1_n_13 ;
  wire \frame_64_transed_reg[0]_i_1_n_14 ;
  wire \frame_64_transed_reg[0]_i_1_n_15 ;
  wire \frame_64_transed_reg[0]_i_1_n_2 ;
  wire \frame_64_transed_reg[0]_i_1_n_3 ;
  wire \frame_64_transed_reg[0]_i_1_n_4 ;
  wire \frame_64_transed_reg[0]_i_1_n_5 ;
  wire \frame_64_transed_reg[0]_i_1_n_6 ;
  wire \frame_64_transed_reg[0]_i_1_n_7 ;
  wire \frame_64_transed_reg[0]_i_1_n_8 ;
  wire \frame_64_transed_reg[0]_i_1_n_9 ;
  wire \frame_64_transed_reg[16]_i_1_n_0 ;
  wire \frame_64_transed_reg[16]_i_1_n_1 ;
  wire \frame_64_transed_reg[16]_i_1_n_10 ;
  wire \frame_64_transed_reg[16]_i_1_n_11 ;
  wire \frame_64_transed_reg[16]_i_1_n_12 ;
  wire \frame_64_transed_reg[16]_i_1_n_13 ;
  wire \frame_64_transed_reg[16]_i_1_n_14 ;
  wire \frame_64_transed_reg[16]_i_1_n_15 ;
  wire \frame_64_transed_reg[16]_i_1_n_2 ;
  wire \frame_64_transed_reg[16]_i_1_n_3 ;
  wire \frame_64_transed_reg[16]_i_1_n_4 ;
  wire \frame_64_transed_reg[16]_i_1_n_5 ;
  wire \frame_64_transed_reg[16]_i_1_n_6 ;
  wire \frame_64_transed_reg[16]_i_1_n_7 ;
  wire \frame_64_transed_reg[16]_i_1_n_8 ;
  wire \frame_64_transed_reg[16]_i_1_n_9 ;
  wire \frame_64_transed_reg[24]_i_1_n_0 ;
  wire \frame_64_transed_reg[24]_i_1_n_1 ;
  wire \frame_64_transed_reg[24]_i_1_n_10 ;
  wire \frame_64_transed_reg[24]_i_1_n_11 ;
  wire \frame_64_transed_reg[24]_i_1_n_12 ;
  wire \frame_64_transed_reg[24]_i_1_n_13 ;
  wire \frame_64_transed_reg[24]_i_1_n_14 ;
  wire \frame_64_transed_reg[24]_i_1_n_15 ;
  wire \frame_64_transed_reg[24]_i_1_n_2 ;
  wire \frame_64_transed_reg[24]_i_1_n_3 ;
  wire \frame_64_transed_reg[24]_i_1_n_4 ;
  wire \frame_64_transed_reg[24]_i_1_n_5 ;
  wire \frame_64_transed_reg[24]_i_1_n_6 ;
  wire \frame_64_transed_reg[24]_i_1_n_7 ;
  wire \frame_64_transed_reg[24]_i_1_n_8 ;
  wire \frame_64_transed_reg[24]_i_1_n_9 ;
  wire \frame_64_transed_reg[32]_i_1_n_0 ;
  wire \frame_64_transed_reg[32]_i_1_n_1 ;
  wire \frame_64_transed_reg[32]_i_1_n_10 ;
  wire \frame_64_transed_reg[32]_i_1_n_11 ;
  wire \frame_64_transed_reg[32]_i_1_n_12 ;
  wire \frame_64_transed_reg[32]_i_1_n_13 ;
  wire \frame_64_transed_reg[32]_i_1_n_14 ;
  wire \frame_64_transed_reg[32]_i_1_n_15 ;
  wire \frame_64_transed_reg[32]_i_1_n_2 ;
  wire \frame_64_transed_reg[32]_i_1_n_3 ;
  wire \frame_64_transed_reg[32]_i_1_n_4 ;
  wire \frame_64_transed_reg[32]_i_1_n_5 ;
  wire \frame_64_transed_reg[32]_i_1_n_6 ;
  wire \frame_64_transed_reg[32]_i_1_n_7 ;
  wire \frame_64_transed_reg[32]_i_1_n_8 ;
  wire \frame_64_transed_reg[32]_i_1_n_9 ;
  wire \frame_64_transed_reg[40]_i_1_n_0 ;
  wire \frame_64_transed_reg[40]_i_1_n_1 ;
  wire \frame_64_transed_reg[40]_i_1_n_10 ;
  wire \frame_64_transed_reg[40]_i_1_n_11 ;
  wire \frame_64_transed_reg[40]_i_1_n_12 ;
  wire \frame_64_transed_reg[40]_i_1_n_13 ;
  wire \frame_64_transed_reg[40]_i_1_n_14 ;
  wire \frame_64_transed_reg[40]_i_1_n_15 ;
  wire \frame_64_transed_reg[40]_i_1_n_2 ;
  wire \frame_64_transed_reg[40]_i_1_n_3 ;
  wire \frame_64_transed_reg[40]_i_1_n_4 ;
  wire \frame_64_transed_reg[40]_i_1_n_5 ;
  wire \frame_64_transed_reg[40]_i_1_n_6 ;
  wire \frame_64_transed_reg[40]_i_1_n_7 ;
  wire \frame_64_transed_reg[40]_i_1_n_8 ;
  wire \frame_64_transed_reg[40]_i_1_n_9 ;
  wire \frame_64_transed_reg[48]_i_1_n_0 ;
  wire \frame_64_transed_reg[48]_i_1_n_1 ;
  wire \frame_64_transed_reg[48]_i_1_n_10 ;
  wire \frame_64_transed_reg[48]_i_1_n_11 ;
  wire \frame_64_transed_reg[48]_i_1_n_12 ;
  wire \frame_64_transed_reg[48]_i_1_n_13 ;
  wire \frame_64_transed_reg[48]_i_1_n_14 ;
  wire \frame_64_transed_reg[48]_i_1_n_15 ;
  wire \frame_64_transed_reg[48]_i_1_n_2 ;
  wire \frame_64_transed_reg[48]_i_1_n_3 ;
  wire \frame_64_transed_reg[48]_i_1_n_4 ;
  wire \frame_64_transed_reg[48]_i_1_n_5 ;
  wire \frame_64_transed_reg[48]_i_1_n_6 ;
  wire \frame_64_transed_reg[48]_i_1_n_7 ;
  wire \frame_64_transed_reg[48]_i_1_n_8 ;
  wire \frame_64_transed_reg[48]_i_1_n_9 ;
  wire \frame_64_transed_reg[56]_i_1_n_1 ;
  wire \frame_64_transed_reg[56]_i_1_n_10 ;
  wire \frame_64_transed_reg[56]_i_1_n_11 ;
  wire \frame_64_transed_reg[56]_i_1_n_12 ;
  wire \frame_64_transed_reg[56]_i_1_n_13 ;
  wire \frame_64_transed_reg[56]_i_1_n_14 ;
  wire \frame_64_transed_reg[56]_i_1_n_15 ;
  wire \frame_64_transed_reg[56]_i_1_n_2 ;
  wire \frame_64_transed_reg[56]_i_1_n_3 ;
  wire \frame_64_transed_reg[56]_i_1_n_4 ;
  wire \frame_64_transed_reg[56]_i_1_n_5 ;
  wire \frame_64_transed_reg[56]_i_1_n_6 ;
  wire \frame_64_transed_reg[56]_i_1_n_7 ;
  wire \frame_64_transed_reg[56]_i_1_n_8 ;
  wire \frame_64_transed_reg[56]_i_1_n_9 ;
  wire \frame_64_transed_reg[8]_i_1_n_0 ;
  wire \frame_64_transed_reg[8]_i_1_n_1 ;
  wire \frame_64_transed_reg[8]_i_1_n_10 ;
  wire \frame_64_transed_reg[8]_i_1_n_11 ;
  wire \frame_64_transed_reg[8]_i_1_n_12 ;
  wire \frame_64_transed_reg[8]_i_1_n_13 ;
  wire \frame_64_transed_reg[8]_i_1_n_14 ;
  wire \frame_64_transed_reg[8]_i_1_n_15 ;
  wire \frame_64_transed_reg[8]_i_1_n_2 ;
  wire \frame_64_transed_reg[8]_i_1_n_3 ;
  wire \frame_64_transed_reg[8]_i_1_n_4 ;
  wire \frame_64_transed_reg[8]_i_1_n_5 ;
  wire \frame_64_transed_reg[8]_i_1_n_6 ;
  wire \frame_64_transed_reg[8]_i_1_n_7 ;
  wire \frame_64_transed_reg[8]_i_1_n_8 ;
  wire \frame_64_transed_reg[8]_i_1_n_9 ;
  wire \frame_65_127_good[0]_i_2_n_0 ;
  wire [63:0]frame_65_127_good_reg;
  wire \frame_65_127_good_reg[0]_i_1_n_0 ;
  wire \frame_65_127_good_reg[0]_i_1_n_1 ;
  wire \frame_65_127_good_reg[0]_i_1_n_10 ;
  wire \frame_65_127_good_reg[0]_i_1_n_11 ;
  wire \frame_65_127_good_reg[0]_i_1_n_12 ;
  wire \frame_65_127_good_reg[0]_i_1_n_13 ;
  wire \frame_65_127_good_reg[0]_i_1_n_14 ;
  wire \frame_65_127_good_reg[0]_i_1_n_15 ;
  wire \frame_65_127_good_reg[0]_i_1_n_2 ;
  wire \frame_65_127_good_reg[0]_i_1_n_3 ;
  wire \frame_65_127_good_reg[0]_i_1_n_4 ;
  wire \frame_65_127_good_reg[0]_i_1_n_5 ;
  wire \frame_65_127_good_reg[0]_i_1_n_6 ;
  wire \frame_65_127_good_reg[0]_i_1_n_7 ;
  wire \frame_65_127_good_reg[0]_i_1_n_8 ;
  wire \frame_65_127_good_reg[0]_i_1_n_9 ;
  wire \frame_65_127_good_reg[16]_i_1_n_0 ;
  wire \frame_65_127_good_reg[16]_i_1_n_1 ;
  wire \frame_65_127_good_reg[16]_i_1_n_10 ;
  wire \frame_65_127_good_reg[16]_i_1_n_11 ;
  wire \frame_65_127_good_reg[16]_i_1_n_12 ;
  wire \frame_65_127_good_reg[16]_i_1_n_13 ;
  wire \frame_65_127_good_reg[16]_i_1_n_14 ;
  wire \frame_65_127_good_reg[16]_i_1_n_15 ;
  wire \frame_65_127_good_reg[16]_i_1_n_2 ;
  wire \frame_65_127_good_reg[16]_i_1_n_3 ;
  wire \frame_65_127_good_reg[16]_i_1_n_4 ;
  wire \frame_65_127_good_reg[16]_i_1_n_5 ;
  wire \frame_65_127_good_reg[16]_i_1_n_6 ;
  wire \frame_65_127_good_reg[16]_i_1_n_7 ;
  wire \frame_65_127_good_reg[16]_i_1_n_8 ;
  wire \frame_65_127_good_reg[16]_i_1_n_9 ;
  wire \frame_65_127_good_reg[24]_i_1_n_0 ;
  wire \frame_65_127_good_reg[24]_i_1_n_1 ;
  wire \frame_65_127_good_reg[24]_i_1_n_10 ;
  wire \frame_65_127_good_reg[24]_i_1_n_11 ;
  wire \frame_65_127_good_reg[24]_i_1_n_12 ;
  wire \frame_65_127_good_reg[24]_i_1_n_13 ;
  wire \frame_65_127_good_reg[24]_i_1_n_14 ;
  wire \frame_65_127_good_reg[24]_i_1_n_15 ;
  wire \frame_65_127_good_reg[24]_i_1_n_2 ;
  wire \frame_65_127_good_reg[24]_i_1_n_3 ;
  wire \frame_65_127_good_reg[24]_i_1_n_4 ;
  wire \frame_65_127_good_reg[24]_i_1_n_5 ;
  wire \frame_65_127_good_reg[24]_i_1_n_6 ;
  wire \frame_65_127_good_reg[24]_i_1_n_7 ;
  wire \frame_65_127_good_reg[24]_i_1_n_8 ;
  wire \frame_65_127_good_reg[24]_i_1_n_9 ;
  wire \frame_65_127_good_reg[32]_i_1_n_0 ;
  wire \frame_65_127_good_reg[32]_i_1_n_1 ;
  wire \frame_65_127_good_reg[32]_i_1_n_10 ;
  wire \frame_65_127_good_reg[32]_i_1_n_11 ;
  wire \frame_65_127_good_reg[32]_i_1_n_12 ;
  wire \frame_65_127_good_reg[32]_i_1_n_13 ;
  wire \frame_65_127_good_reg[32]_i_1_n_14 ;
  wire \frame_65_127_good_reg[32]_i_1_n_15 ;
  wire \frame_65_127_good_reg[32]_i_1_n_2 ;
  wire \frame_65_127_good_reg[32]_i_1_n_3 ;
  wire \frame_65_127_good_reg[32]_i_1_n_4 ;
  wire \frame_65_127_good_reg[32]_i_1_n_5 ;
  wire \frame_65_127_good_reg[32]_i_1_n_6 ;
  wire \frame_65_127_good_reg[32]_i_1_n_7 ;
  wire \frame_65_127_good_reg[32]_i_1_n_8 ;
  wire \frame_65_127_good_reg[32]_i_1_n_9 ;
  wire \frame_65_127_good_reg[40]_i_1_n_0 ;
  wire \frame_65_127_good_reg[40]_i_1_n_1 ;
  wire \frame_65_127_good_reg[40]_i_1_n_10 ;
  wire \frame_65_127_good_reg[40]_i_1_n_11 ;
  wire \frame_65_127_good_reg[40]_i_1_n_12 ;
  wire \frame_65_127_good_reg[40]_i_1_n_13 ;
  wire \frame_65_127_good_reg[40]_i_1_n_14 ;
  wire \frame_65_127_good_reg[40]_i_1_n_15 ;
  wire \frame_65_127_good_reg[40]_i_1_n_2 ;
  wire \frame_65_127_good_reg[40]_i_1_n_3 ;
  wire \frame_65_127_good_reg[40]_i_1_n_4 ;
  wire \frame_65_127_good_reg[40]_i_1_n_5 ;
  wire \frame_65_127_good_reg[40]_i_1_n_6 ;
  wire \frame_65_127_good_reg[40]_i_1_n_7 ;
  wire \frame_65_127_good_reg[40]_i_1_n_8 ;
  wire \frame_65_127_good_reg[40]_i_1_n_9 ;
  wire \frame_65_127_good_reg[48]_i_1_n_0 ;
  wire \frame_65_127_good_reg[48]_i_1_n_1 ;
  wire \frame_65_127_good_reg[48]_i_1_n_10 ;
  wire \frame_65_127_good_reg[48]_i_1_n_11 ;
  wire \frame_65_127_good_reg[48]_i_1_n_12 ;
  wire \frame_65_127_good_reg[48]_i_1_n_13 ;
  wire \frame_65_127_good_reg[48]_i_1_n_14 ;
  wire \frame_65_127_good_reg[48]_i_1_n_15 ;
  wire \frame_65_127_good_reg[48]_i_1_n_2 ;
  wire \frame_65_127_good_reg[48]_i_1_n_3 ;
  wire \frame_65_127_good_reg[48]_i_1_n_4 ;
  wire \frame_65_127_good_reg[48]_i_1_n_5 ;
  wire \frame_65_127_good_reg[48]_i_1_n_6 ;
  wire \frame_65_127_good_reg[48]_i_1_n_7 ;
  wire \frame_65_127_good_reg[48]_i_1_n_8 ;
  wire \frame_65_127_good_reg[48]_i_1_n_9 ;
  wire \frame_65_127_good_reg[56]_i_1_n_1 ;
  wire \frame_65_127_good_reg[56]_i_1_n_10 ;
  wire \frame_65_127_good_reg[56]_i_1_n_11 ;
  wire \frame_65_127_good_reg[56]_i_1_n_12 ;
  wire \frame_65_127_good_reg[56]_i_1_n_13 ;
  wire \frame_65_127_good_reg[56]_i_1_n_14 ;
  wire \frame_65_127_good_reg[56]_i_1_n_15 ;
  wire \frame_65_127_good_reg[56]_i_1_n_2 ;
  wire \frame_65_127_good_reg[56]_i_1_n_3 ;
  wire \frame_65_127_good_reg[56]_i_1_n_4 ;
  wire \frame_65_127_good_reg[56]_i_1_n_5 ;
  wire \frame_65_127_good_reg[56]_i_1_n_6 ;
  wire \frame_65_127_good_reg[56]_i_1_n_7 ;
  wire \frame_65_127_good_reg[56]_i_1_n_8 ;
  wire \frame_65_127_good_reg[56]_i_1_n_9 ;
  wire \frame_65_127_good_reg[8]_i_1_n_0 ;
  wire \frame_65_127_good_reg[8]_i_1_n_1 ;
  wire \frame_65_127_good_reg[8]_i_1_n_10 ;
  wire \frame_65_127_good_reg[8]_i_1_n_11 ;
  wire \frame_65_127_good_reg[8]_i_1_n_12 ;
  wire \frame_65_127_good_reg[8]_i_1_n_13 ;
  wire \frame_65_127_good_reg[8]_i_1_n_14 ;
  wire \frame_65_127_good_reg[8]_i_1_n_15 ;
  wire \frame_65_127_good_reg[8]_i_1_n_2 ;
  wire \frame_65_127_good_reg[8]_i_1_n_3 ;
  wire \frame_65_127_good_reg[8]_i_1_n_4 ;
  wire \frame_65_127_good_reg[8]_i_1_n_5 ;
  wire \frame_65_127_good_reg[8]_i_1_n_6 ;
  wire \frame_65_127_good_reg[8]_i_1_n_7 ;
  wire \frame_65_127_good_reg[8]_i_1_n_8 ;
  wire \frame_65_127_good_reg[8]_i_1_n_9 ;
  wire \frame_65_127_transed[0]_i_2_n_0 ;
  wire [63:0]frame_65_127_transed_reg;
  wire \frame_65_127_transed_reg[0]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[0]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[16]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[24]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[32]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[40]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[48]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[56]_i_1_n_9 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_0 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_1 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_10 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_11 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_12 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_13 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_14 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_15 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_2 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_3 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_4 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_5 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_6 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_7 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_8 ;
  wire \frame_65_127_transed_reg[8]_i_1_n_9 ;
  wire \frame_received_good[0]_i_2_n_0 ;
  wire [63:0]frame_received_good_reg;
  wire \frame_received_good_reg[0]_i_1_n_0 ;
  wire \frame_received_good_reg[0]_i_1_n_1 ;
  wire \frame_received_good_reg[0]_i_1_n_10 ;
  wire \frame_received_good_reg[0]_i_1_n_11 ;
  wire \frame_received_good_reg[0]_i_1_n_12 ;
  wire \frame_received_good_reg[0]_i_1_n_13 ;
  wire \frame_received_good_reg[0]_i_1_n_14 ;
  wire \frame_received_good_reg[0]_i_1_n_15 ;
  wire \frame_received_good_reg[0]_i_1_n_2 ;
  wire \frame_received_good_reg[0]_i_1_n_3 ;
  wire \frame_received_good_reg[0]_i_1_n_4 ;
  wire \frame_received_good_reg[0]_i_1_n_5 ;
  wire \frame_received_good_reg[0]_i_1_n_6 ;
  wire \frame_received_good_reg[0]_i_1_n_7 ;
  wire \frame_received_good_reg[0]_i_1_n_8 ;
  wire \frame_received_good_reg[0]_i_1_n_9 ;
  wire \frame_received_good_reg[16]_i_1_n_0 ;
  wire \frame_received_good_reg[16]_i_1_n_1 ;
  wire \frame_received_good_reg[16]_i_1_n_10 ;
  wire \frame_received_good_reg[16]_i_1_n_11 ;
  wire \frame_received_good_reg[16]_i_1_n_12 ;
  wire \frame_received_good_reg[16]_i_1_n_13 ;
  wire \frame_received_good_reg[16]_i_1_n_14 ;
  wire \frame_received_good_reg[16]_i_1_n_15 ;
  wire \frame_received_good_reg[16]_i_1_n_2 ;
  wire \frame_received_good_reg[16]_i_1_n_3 ;
  wire \frame_received_good_reg[16]_i_1_n_4 ;
  wire \frame_received_good_reg[16]_i_1_n_5 ;
  wire \frame_received_good_reg[16]_i_1_n_6 ;
  wire \frame_received_good_reg[16]_i_1_n_7 ;
  wire \frame_received_good_reg[16]_i_1_n_8 ;
  wire \frame_received_good_reg[16]_i_1_n_9 ;
  wire \frame_received_good_reg[24]_i_1_n_0 ;
  wire \frame_received_good_reg[24]_i_1_n_1 ;
  wire \frame_received_good_reg[24]_i_1_n_10 ;
  wire \frame_received_good_reg[24]_i_1_n_11 ;
  wire \frame_received_good_reg[24]_i_1_n_12 ;
  wire \frame_received_good_reg[24]_i_1_n_13 ;
  wire \frame_received_good_reg[24]_i_1_n_14 ;
  wire \frame_received_good_reg[24]_i_1_n_15 ;
  wire \frame_received_good_reg[24]_i_1_n_2 ;
  wire \frame_received_good_reg[24]_i_1_n_3 ;
  wire \frame_received_good_reg[24]_i_1_n_4 ;
  wire \frame_received_good_reg[24]_i_1_n_5 ;
  wire \frame_received_good_reg[24]_i_1_n_6 ;
  wire \frame_received_good_reg[24]_i_1_n_7 ;
  wire \frame_received_good_reg[24]_i_1_n_8 ;
  wire \frame_received_good_reg[24]_i_1_n_9 ;
  wire \frame_received_good_reg[32]_i_1_n_0 ;
  wire \frame_received_good_reg[32]_i_1_n_1 ;
  wire \frame_received_good_reg[32]_i_1_n_10 ;
  wire \frame_received_good_reg[32]_i_1_n_11 ;
  wire \frame_received_good_reg[32]_i_1_n_12 ;
  wire \frame_received_good_reg[32]_i_1_n_13 ;
  wire \frame_received_good_reg[32]_i_1_n_14 ;
  wire \frame_received_good_reg[32]_i_1_n_15 ;
  wire \frame_received_good_reg[32]_i_1_n_2 ;
  wire \frame_received_good_reg[32]_i_1_n_3 ;
  wire \frame_received_good_reg[32]_i_1_n_4 ;
  wire \frame_received_good_reg[32]_i_1_n_5 ;
  wire \frame_received_good_reg[32]_i_1_n_6 ;
  wire \frame_received_good_reg[32]_i_1_n_7 ;
  wire \frame_received_good_reg[32]_i_1_n_8 ;
  wire \frame_received_good_reg[32]_i_1_n_9 ;
  wire \frame_received_good_reg[40]_i_1_n_0 ;
  wire \frame_received_good_reg[40]_i_1_n_1 ;
  wire \frame_received_good_reg[40]_i_1_n_10 ;
  wire \frame_received_good_reg[40]_i_1_n_11 ;
  wire \frame_received_good_reg[40]_i_1_n_12 ;
  wire \frame_received_good_reg[40]_i_1_n_13 ;
  wire \frame_received_good_reg[40]_i_1_n_14 ;
  wire \frame_received_good_reg[40]_i_1_n_15 ;
  wire \frame_received_good_reg[40]_i_1_n_2 ;
  wire \frame_received_good_reg[40]_i_1_n_3 ;
  wire \frame_received_good_reg[40]_i_1_n_4 ;
  wire \frame_received_good_reg[40]_i_1_n_5 ;
  wire \frame_received_good_reg[40]_i_1_n_6 ;
  wire \frame_received_good_reg[40]_i_1_n_7 ;
  wire \frame_received_good_reg[40]_i_1_n_8 ;
  wire \frame_received_good_reg[40]_i_1_n_9 ;
  wire \frame_received_good_reg[48]_i_1_n_0 ;
  wire \frame_received_good_reg[48]_i_1_n_1 ;
  wire \frame_received_good_reg[48]_i_1_n_10 ;
  wire \frame_received_good_reg[48]_i_1_n_11 ;
  wire \frame_received_good_reg[48]_i_1_n_12 ;
  wire \frame_received_good_reg[48]_i_1_n_13 ;
  wire \frame_received_good_reg[48]_i_1_n_14 ;
  wire \frame_received_good_reg[48]_i_1_n_15 ;
  wire \frame_received_good_reg[48]_i_1_n_2 ;
  wire \frame_received_good_reg[48]_i_1_n_3 ;
  wire \frame_received_good_reg[48]_i_1_n_4 ;
  wire \frame_received_good_reg[48]_i_1_n_5 ;
  wire \frame_received_good_reg[48]_i_1_n_6 ;
  wire \frame_received_good_reg[48]_i_1_n_7 ;
  wire \frame_received_good_reg[48]_i_1_n_8 ;
  wire \frame_received_good_reg[48]_i_1_n_9 ;
  wire \frame_received_good_reg[56]_i_1_n_1 ;
  wire \frame_received_good_reg[56]_i_1_n_10 ;
  wire \frame_received_good_reg[56]_i_1_n_11 ;
  wire \frame_received_good_reg[56]_i_1_n_12 ;
  wire \frame_received_good_reg[56]_i_1_n_13 ;
  wire \frame_received_good_reg[56]_i_1_n_14 ;
  wire \frame_received_good_reg[56]_i_1_n_15 ;
  wire \frame_received_good_reg[56]_i_1_n_2 ;
  wire \frame_received_good_reg[56]_i_1_n_3 ;
  wire \frame_received_good_reg[56]_i_1_n_4 ;
  wire \frame_received_good_reg[56]_i_1_n_5 ;
  wire \frame_received_good_reg[56]_i_1_n_6 ;
  wire \frame_received_good_reg[56]_i_1_n_7 ;
  wire \frame_received_good_reg[56]_i_1_n_8 ;
  wire \frame_received_good_reg[56]_i_1_n_9 ;
  wire \frame_received_good_reg[8]_i_1_n_0 ;
  wire \frame_received_good_reg[8]_i_1_n_1 ;
  wire \frame_received_good_reg[8]_i_1_n_10 ;
  wire \frame_received_good_reg[8]_i_1_n_11 ;
  wire \frame_received_good_reg[8]_i_1_n_12 ;
  wire \frame_received_good_reg[8]_i_1_n_13 ;
  wire \frame_received_good_reg[8]_i_1_n_14 ;
  wire \frame_received_good_reg[8]_i_1_n_15 ;
  wire \frame_received_good_reg[8]_i_1_n_2 ;
  wire \frame_received_good_reg[8]_i_1_n_3 ;
  wire \frame_received_good_reg[8]_i_1_n_4 ;
  wire \frame_received_good_reg[8]_i_1_n_5 ;
  wire \frame_received_good_reg[8]_i_1_n_6 ;
  wire \frame_received_good_reg[8]_i_1_n_7 ;
  wire \frame_received_good_reg[8]_i_1_n_8 ;
  wire \frame_received_good_reg[8]_i_1_n_9 ;
  wire \good_frame_transed[0]_i_2_n_0 ;
  wire [63:0]good_frame_transed_reg;
  wire \good_frame_transed_reg[0]_i_1_n_0 ;
  wire \good_frame_transed_reg[0]_i_1_n_1 ;
  wire \good_frame_transed_reg[0]_i_1_n_10 ;
  wire \good_frame_transed_reg[0]_i_1_n_11 ;
  wire \good_frame_transed_reg[0]_i_1_n_12 ;
  wire \good_frame_transed_reg[0]_i_1_n_13 ;
  wire \good_frame_transed_reg[0]_i_1_n_14 ;
  wire \good_frame_transed_reg[0]_i_1_n_15 ;
  wire \good_frame_transed_reg[0]_i_1_n_2 ;
  wire \good_frame_transed_reg[0]_i_1_n_3 ;
  wire \good_frame_transed_reg[0]_i_1_n_4 ;
  wire \good_frame_transed_reg[0]_i_1_n_5 ;
  wire \good_frame_transed_reg[0]_i_1_n_6 ;
  wire \good_frame_transed_reg[0]_i_1_n_7 ;
  wire \good_frame_transed_reg[0]_i_1_n_8 ;
  wire \good_frame_transed_reg[0]_i_1_n_9 ;
  wire \good_frame_transed_reg[16]_i_1_n_0 ;
  wire \good_frame_transed_reg[16]_i_1_n_1 ;
  wire \good_frame_transed_reg[16]_i_1_n_10 ;
  wire \good_frame_transed_reg[16]_i_1_n_11 ;
  wire \good_frame_transed_reg[16]_i_1_n_12 ;
  wire \good_frame_transed_reg[16]_i_1_n_13 ;
  wire \good_frame_transed_reg[16]_i_1_n_14 ;
  wire \good_frame_transed_reg[16]_i_1_n_15 ;
  wire \good_frame_transed_reg[16]_i_1_n_2 ;
  wire \good_frame_transed_reg[16]_i_1_n_3 ;
  wire \good_frame_transed_reg[16]_i_1_n_4 ;
  wire \good_frame_transed_reg[16]_i_1_n_5 ;
  wire \good_frame_transed_reg[16]_i_1_n_6 ;
  wire \good_frame_transed_reg[16]_i_1_n_7 ;
  wire \good_frame_transed_reg[16]_i_1_n_8 ;
  wire \good_frame_transed_reg[16]_i_1_n_9 ;
  wire \good_frame_transed_reg[24]_i_1_n_0 ;
  wire \good_frame_transed_reg[24]_i_1_n_1 ;
  wire \good_frame_transed_reg[24]_i_1_n_10 ;
  wire \good_frame_transed_reg[24]_i_1_n_11 ;
  wire \good_frame_transed_reg[24]_i_1_n_12 ;
  wire \good_frame_transed_reg[24]_i_1_n_13 ;
  wire \good_frame_transed_reg[24]_i_1_n_14 ;
  wire \good_frame_transed_reg[24]_i_1_n_15 ;
  wire \good_frame_transed_reg[24]_i_1_n_2 ;
  wire \good_frame_transed_reg[24]_i_1_n_3 ;
  wire \good_frame_transed_reg[24]_i_1_n_4 ;
  wire \good_frame_transed_reg[24]_i_1_n_5 ;
  wire \good_frame_transed_reg[24]_i_1_n_6 ;
  wire \good_frame_transed_reg[24]_i_1_n_7 ;
  wire \good_frame_transed_reg[24]_i_1_n_8 ;
  wire \good_frame_transed_reg[24]_i_1_n_9 ;
  wire \good_frame_transed_reg[32]_i_1_n_0 ;
  wire \good_frame_transed_reg[32]_i_1_n_1 ;
  wire \good_frame_transed_reg[32]_i_1_n_10 ;
  wire \good_frame_transed_reg[32]_i_1_n_11 ;
  wire \good_frame_transed_reg[32]_i_1_n_12 ;
  wire \good_frame_transed_reg[32]_i_1_n_13 ;
  wire \good_frame_transed_reg[32]_i_1_n_14 ;
  wire \good_frame_transed_reg[32]_i_1_n_15 ;
  wire \good_frame_transed_reg[32]_i_1_n_2 ;
  wire \good_frame_transed_reg[32]_i_1_n_3 ;
  wire \good_frame_transed_reg[32]_i_1_n_4 ;
  wire \good_frame_transed_reg[32]_i_1_n_5 ;
  wire \good_frame_transed_reg[32]_i_1_n_6 ;
  wire \good_frame_transed_reg[32]_i_1_n_7 ;
  wire \good_frame_transed_reg[32]_i_1_n_8 ;
  wire \good_frame_transed_reg[32]_i_1_n_9 ;
  wire \good_frame_transed_reg[40]_i_1_n_0 ;
  wire \good_frame_transed_reg[40]_i_1_n_1 ;
  wire \good_frame_transed_reg[40]_i_1_n_10 ;
  wire \good_frame_transed_reg[40]_i_1_n_11 ;
  wire \good_frame_transed_reg[40]_i_1_n_12 ;
  wire \good_frame_transed_reg[40]_i_1_n_13 ;
  wire \good_frame_transed_reg[40]_i_1_n_14 ;
  wire \good_frame_transed_reg[40]_i_1_n_15 ;
  wire \good_frame_transed_reg[40]_i_1_n_2 ;
  wire \good_frame_transed_reg[40]_i_1_n_3 ;
  wire \good_frame_transed_reg[40]_i_1_n_4 ;
  wire \good_frame_transed_reg[40]_i_1_n_5 ;
  wire \good_frame_transed_reg[40]_i_1_n_6 ;
  wire \good_frame_transed_reg[40]_i_1_n_7 ;
  wire \good_frame_transed_reg[40]_i_1_n_8 ;
  wire \good_frame_transed_reg[40]_i_1_n_9 ;
  wire \good_frame_transed_reg[48]_i_1_n_0 ;
  wire \good_frame_transed_reg[48]_i_1_n_1 ;
  wire \good_frame_transed_reg[48]_i_1_n_10 ;
  wire \good_frame_transed_reg[48]_i_1_n_11 ;
  wire \good_frame_transed_reg[48]_i_1_n_12 ;
  wire \good_frame_transed_reg[48]_i_1_n_13 ;
  wire \good_frame_transed_reg[48]_i_1_n_14 ;
  wire \good_frame_transed_reg[48]_i_1_n_15 ;
  wire \good_frame_transed_reg[48]_i_1_n_2 ;
  wire \good_frame_transed_reg[48]_i_1_n_3 ;
  wire \good_frame_transed_reg[48]_i_1_n_4 ;
  wire \good_frame_transed_reg[48]_i_1_n_5 ;
  wire \good_frame_transed_reg[48]_i_1_n_6 ;
  wire \good_frame_transed_reg[48]_i_1_n_7 ;
  wire \good_frame_transed_reg[48]_i_1_n_8 ;
  wire \good_frame_transed_reg[48]_i_1_n_9 ;
  wire \good_frame_transed_reg[56]_i_1_n_1 ;
  wire \good_frame_transed_reg[56]_i_1_n_10 ;
  wire \good_frame_transed_reg[56]_i_1_n_11 ;
  wire \good_frame_transed_reg[56]_i_1_n_12 ;
  wire \good_frame_transed_reg[56]_i_1_n_13 ;
  wire \good_frame_transed_reg[56]_i_1_n_14 ;
  wire \good_frame_transed_reg[56]_i_1_n_15 ;
  wire \good_frame_transed_reg[56]_i_1_n_2 ;
  wire \good_frame_transed_reg[56]_i_1_n_3 ;
  wire \good_frame_transed_reg[56]_i_1_n_4 ;
  wire \good_frame_transed_reg[56]_i_1_n_5 ;
  wire \good_frame_transed_reg[56]_i_1_n_6 ;
  wire \good_frame_transed_reg[56]_i_1_n_7 ;
  wire \good_frame_transed_reg[56]_i_1_n_8 ;
  wire \good_frame_transed_reg[56]_i_1_n_9 ;
  wire \good_frame_transed_reg[8]_i_1_n_0 ;
  wire \good_frame_transed_reg[8]_i_1_n_1 ;
  wire \good_frame_transed_reg[8]_i_1_n_10 ;
  wire \good_frame_transed_reg[8]_i_1_n_11 ;
  wire \good_frame_transed_reg[8]_i_1_n_12 ;
  wire \good_frame_transed_reg[8]_i_1_n_13 ;
  wire \good_frame_transed_reg[8]_i_1_n_14 ;
  wire \good_frame_transed_reg[8]_i_1_n_15 ;
  wire \good_frame_transed_reg[8]_i_1_n_2 ;
  wire \good_frame_transed_reg[8]_i_1_n_3 ;
  wire \good_frame_transed_reg[8]_i_1_n_4 ;
  wire \good_frame_transed_reg[8]_i_1_n_5 ;
  wire \good_frame_transed_reg[8]_i_1_n_6 ;
  wire \good_frame_transed_reg[8]_i_1_n_7 ;
  wire \good_frame_transed_reg[8]_i_1_n_8 ;
  wire \good_frame_transed_reg[8]_i_1_n_9 ;
  wire in0;
  wire \lt_out_range[0]_i_2_n_0 ;
  wire [63:0]lt_out_range_reg;
  wire \lt_out_range_reg[0]_i_1_n_0 ;
  wire \lt_out_range_reg[0]_i_1_n_1 ;
  wire \lt_out_range_reg[0]_i_1_n_10 ;
  wire \lt_out_range_reg[0]_i_1_n_11 ;
  wire \lt_out_range_reg[0]_i_1_n_12 ;
  wire \lt_out_range_reg[0]_i_1_n_13 ;
  wire \lt_out_range_reg[0]_i_1_n_14 ;
  wire \lt_out_range_reg[0]_i_1_n_15 ;
  wire \lt_out_range_reg[0]_i_1_n_2 ;
  wire \lt_out_range_reg[0]_i_1_n_3 ;
  wire \lt_out_range_reg[0]_i_1_n_4 ;
  wire \lt_out_range_reg[0]_i_1_n_5 ;
  wire \lt_out_range_reg[0]_i_1_n_6 ;
  wire \lt_out_range_reg[0]_i_1_n_7 ;
  wire \lt_out_range_reg[0]_i_1_n_8 ;
  wire \lt_out_range_reg[0]_i_1_n_9 ;
  wire \lt_out_range_reg[16]_i_1_n_0 ;
  wire \lt_out_range_reg[16]_i_1_n_1 ;
  wire \lt_out_range_reg[16]_i_1_n_10 ;
  wire \lt_out_range_reg[16]_i_1_n_11 ;
  wire \lt_out_range_reg[16]_i_1_n_12 ;
  wire \lt_out_range_reg[16]_i_1_n_13 ;
  wire \lt_out_range_reg[16]_i_1_n_14 ;
  wire \lt_out_range_reg[16]_i_1_n_15 ;
  wire \lt_out_range_reg[16]_i_1_n_2 ;
  wire \lt_out_range_reg[16]_i_1_n_3 ;
  wire \lt_out_range_reg[16]_i_1_n_4 ;
  wire \lt_out_range_reg[16]_i_1_n_5 ;
  wire \lt_out_range_reg[16]_i_1_n_6 ;
  wire \lt_out_range_reg[16]_i_1_n_7 ;
  wire \lt_out_range_reg[16]_i_1_n_8 ;
  wire \lt_out_range_reg[16]_i_1_n_9 ;
  wire \lt_out_range_reg[24]_i_1_n_0 ;
  wire \lt_out_range_reg[24]_i_1_n_1 ;
  wire \lt_out_range_reg[24]_i_1_n_10 ;
  wire \lt_out_range_reg[24]_i_1_n_11 ;
  wire \lt_out_range_reg[24]_i_1_n_12 ;
  wire \lt_out_range_reg[24]_i_1_n_13 ;
  wire \lt_out_range_reg[24]_i_1_n_14 ;
  wire \lt_out_range_reg[24]_i_1_n_15 ;
  wire \lt_out_range_reg[24]_i_1_n_2 ;
  wire \lt_out_range_reg[24]_i_1_n_3 ;
  wire \lt_out_range_reg[24]_i_1_n_4 ;
  wire \lt_out_range_reg[24]_i_1_n_5 ;
  wire \lt_out_range_reg[24]_i_1_n_6 ;
  wire \lt_out_range_reg[24]_i_1_n_7 ;
  wire \lt_out_range_reg[24]_i_1_n_8 ;
  wire \lt_out_range_reg[24]_i_1_n_9 ;
  wire \lt_out_range_reg[32]_i_1_n_0 ;
  wire \lt_out_range_reg[32]_i_1_n_1 ;
  wire \lt_out_range_reg[32]_i_1_n_10 ;
  wire \lt_out_range_reg[32]_i_1_n_11 ;
  wire \lt_out_range_reg[32]_i_1_n_12 ;
  wire \lt_out_range_reg[32]_i_1_n_13 ;
  wire \lt_out_range_reg[32]_i_1_n_14 ;
  wire \lt_out_range_reg[32]_i_1_n_15 ;
  wire \lt_out_range_reg[32]_i_1_n_2 ;
  wire \lt_out_range_reg[32]_i_1_n_3 ;
  wire \lt_out_range_reg[32]_i_1_n_4 ;
  wire \lt_out_range_reg[32]_i_1_n_5 ;
  wire \lt_out_range_reg[32]_i_1_n_6 ;
  wire \lt_out_range_reg[32]_i_1_n_7 ;
  wire \lt_out_range_reg[32]_i_1_n_8 ;
  wire \lt_out_range_reg[32]_i_1_n_9 ;
  wire \lt_out_range_reg[40]_i_1_n_0 ;
  wire \lt_out_range_reg[40]_i_1_n_1 ;
  wire \lt_out_range_reg[40]_i_1_n_10 ;
  wire \lt_out_range_reg[40]_i_1_n_11 ;
  wire \lt_out_range_reg[40]_i_1_n_12 ;
  wire \lt_out_range_reg[40]_i_1_n_13 ;
  wire \lt_out_range_reg[40]_i_1_n_14 ;
  wire \lt_out_range_reg[40]_i_1_n_15 ;
  wire \lt_out_range_reg[40]_i_1_n_2 ;
  wire \lt_out_range_reg[40]_i_1_n_3 ;
  wire \lt_out_range_reg[40]_i_1_n_4 ;
  wire \lt_out_range_reg[40]_i_1_n_5 ;
  wire \lt_out_range_reg[40]_i_1_n_6 ;
  wire \lt_out_range_reg[40]_i_1_n_7 ;
  wire \lt_out_range_reg[40]_i_1_n_8 ;
  wire \lt_out_range_reg[40]_i_1_n_9 ;
  wire \lt_out_range_reg[48]_i_1_n_0 ;
  wire \lt_out_range_reg[48]_i_1_n_1 ;
  wire \lt_out_range_reg[48]_i_1_n_10 ;
  wire \lt_out_range_reg[48]_i_1_n_11 ;
  wire \lt_out_range_reg[48]_i_1_n_12 ;
  wire \lt_out_range_reg[48]_i_1_n_13 ;
  wire \lt_out_range_reg[48]_i_1_n_14 ;
  wire \lt_out_range_reg[48]_i_1_n_15 ;
  wire \lt_out_range_reg[48]_i_1_n_2 ;
  wire \lt_out_range_reg[48]_i_1_n_3 ;
  wire \lt_out_range_reg[48]_i_1_n_4 ;
  wire \lt_out_range_reg[48]_i_1_n_5 ;
  wire \lt_out_range_reg[48]_i_1_n_6 ;
  wire \lt_out_range_reg[48]_i_1_n_7 ;
  wire \lt_out_range_reg[48]_i_1_n_8 ;
  wire \lt_out_range_reg[48]_i_1_n_9 ;
  wire \lt_out_range_reg[56]_i_1_n_1 ;
  wire \lt_out_range_reg[56]_i_1_n_10 ;
  wire \lt_out_range_reg[56]_i_1_n_11 ;
  wire \lt_out_range_reg[56]_i_1_n_12 ;
  wire \lt_out_range_reg[56]_i_1_n_13 ;
  wire \lt_out_range_reg[56]_i_1_n_14 ;
  wire \lt_out_range_reg[56]_i_1_n_15 ;
  wire \lt_out_range_reg[56]_i_1_n_2 ;
  wire \lt_out_range_reg[56]_i_1_n_3 ;
  wire \lt_out_range_reg[56]_i_1_n_4 ;
  wire \lt_out_range_reg[56]_i_1_n_5 ;
  wire \lt_out_range_reg[56]_i_1_n_6 ;
  wire \lt_out_range_reg[56]_i_1_n_7 ;
  wire \lt_out_range_reg[56]_i_1_n_8 ;
  wire \lt_out_range_reg[56]_i_1_n_9 ;
  wire \lt_out_range_reg[8]_i_1_n_0 ;
  wire \lt_out_range_reg[8]_i_1_n_1 ;
  wire \lt_out_range_reg[8]_i_1_n_10 ;
  wire \lt_out_range_reg[8]_i_1_n_11 ;
  wire \lt_out_range_reg[8]_i_1_n_12 ;
  wire \lt_out_range_reg[8]_i_1_n_13 ;
  wire \lt_out_range_reg[8]_i_1_n_14 ;
  wire \lt_out_range_reg[8]_i_1_n_15 ;
  wire \lt_out_range_reg[8]_i_1_n_2 ;
  wire \lt_out_range_reg[8]_i_1_n_3 ;
  wire \lt_out_range_reg[8]_i_1_n_4 ;
  wire \lt_out_range_reg[8]_i_1_n_5 ;
  wire \lt_out_range_reg[8]_i_1_n_6 ;
  wire \lt_out_range_reg[8]_i_1_n_7 ;
  wire \lt_out_range_reg[8]_i_1_n_8 ;
  wire \lt_out_range_reg[8]_i_1_n_9 ;
  wire mdio_in_valid;
  wire mdio_in_valid_d1;
  wire [0:0]mdio_opcode;
  wire \mdio_opcode[1]_i_1_n_0 ;
  wire mdio_out_valid;
  wire mdio_out_valid_i_1_n_0;
  wire mdio_out_valid_i_2_n_0;
  wire [31:5]mgmt_config;
  wire \mgmt_config[31]_i_1_n_0 ;
  wire \mgmt_config[31]_i_2_n_0 ;
  wire mgmt_miim_rdy_i_1_n_0;
  wire [31:0]mgmt_rd_data;
  wire mgmt_rd_data0;
  wire [15:0]mgmt_rd_data0_in;
  wire \mgmt_rd_data[0]_i_2_n_0 ;
  wire \mgmt_rd_data[0]_i_4_n_0 ;
  wire \mgmt_rd_data[10]_i_2_n_0 ;
  wire \mgmt_rd_data[10]_i_4_n_0 ;
  wire \mgmt_rd_data[11]_i_2_n_0 ;
  wire \mgmt_rd_data[11]_i_4_n_0 ;
  wire \mgmt_rd_data[12]_i_2_n_0 ;
  wire \mgmt_rd_data[12]_i_4_n_0 ;
  wire \mgmt_rd_data[13]_i_2_n_0 ;
  wire \mgmt_rd_data[13]_i_4_n_0 ;
  wire \mgmt_rd_data[14]_i_2_n_0 ;
  wire \mgmt_rd_data[14]_i_4_n_0 ;
  wire \mgmt_rd_data[15]_i_2_n_0 ;
  wire \mgmt_rd_data[15]_i_4_n_0 ;
  wire \mgmt_rd_data[16]_i_2_n_0 ;
  wire \mgmt_rd_data[16]_i_3_n_0 ;
  wire \mgmt_rd_data[17]_i_2_n_0 ;
  wire \mgmt_rd_data[17]_i_3_n_0 ;
  wire \mgmt_rd_data[18]_i_2_n_0 ;
  wire \mgmt_rd_data[18]_i_3_n_0 ;
  wire \mgmt_rd_data[19]_i_2_n_0 ;
  wire \mgmt_rd_data[19]_i_3_n_0 ;
  wire \mgmt_rd_data[1]_i_2_n_0 ;
  wire \mgmt_rd_data[1]_i_4_n_0 ;
  wire \mgmt_rd_data[20]_i_2_n_0 ;
  wire \mgmt_rd_data[20]_i_3_n_0 ;
  wire \mgmt_rd_data[21]_i_2_n_0 ;
  wire \mgmt_rd_data[21]_i_3_n_0 ;
  wire \mgmt_rd_data[22]_i_2_n_0 ;
  wire \mgmt_rd_data[22]_i_3_n_0 ;
  wire \mgmt_rd_data[23]_i_2_n_0 ;
  wire \mgmt_rd_data[23]_i_3_n_0 ;
  wire \mgmt_rd_data[24]_i_2_n_0 ;
  wire \mgmt_rd_data[24]_i_3_n_0 ;
  wire \mgmt_rd_data[25]_i_2_n_0 ;
  wire \mgmt_rd_data[25]_i_3_n_0 ;
  wire \mgmt_rd_data[26]_i_2_n_0 ;
  wire \mgmt_rd_data[26]_i_3_n_0 ;
  wire \mgmt_rd_data[27]_i_2_n_0 ;
  wire \mgmt_rd_data[27]_i_3_n_0 ;
  wire \mgmt_rd_data[28]_i_2_n_0 ;
  wire \mgmt_rd_data[28]_i_3_n_0 ;
  wire \mgmt_rd_data[29]_i_2_n_0 ;
  wire \mgmt_rd_data[29]_i_3_n_0 ;
  wire \mgmt_rd_data[2]_i_2_n_0 ;
  wire \mgmt_rd_data[2]_i_4_n_0 ;
  wire \mgmt_rd_data[30]_i_2_n_0 ;
  wire \mgmt_rd_data[30]_i_3_n_0 ;
  wire \mgmt_rd_data[31]_i_3_n_0 ;
  wire \mgmt_rd_data[31]_i_4_n_0 ;
  wire \mgmt_rd_data[31]_i_5_n_0 ;
  wire \mgmt_rd_data[3]_i_2_n_0 ;
  wire \mgmt_rd_data[3]_i_4_n_0 ;
  wire \mgmt_rd_data[4]_i_2_n_0 ;
  wire \mgmt_rd_data[4]_i_4_n_0 ;
  wire \mgmt_rd_data[5]_i_2_n_0 ;
  wire \mgmt_rd_data[5]_i_4_n_0 ;
  wire \mgmt_rd_data[6]_i_2_n_0 ;
  wire \mgmt_rd_data[6]_i_4_n_0 ;
  wire \mgmt_rd_data[7]_i_2_n_0 ;
  wire \mgmt_rd_data[7]_i_4_n_0 ;
  wire \mgmt_rd_data[8]_i_2_n_0 ;
  wire \mgmt_rd_data[8]_i_4_n_0 ;
  wire \mgmt_rd_data[9]_i_2_n_0 ;
  wire \mgmt_rd_data[9]_i_4_n_0 ;
  wire [15:0]\mgmt_rd_data_reg[15]_0 ;
  wire [31:0]mgmt_wr_data;
  wire \multicast_frame_transed[0]_i_2_n_0 ;
  wire [63:0]multicast_frame_transed_reg;
  wire \multicast_frame_transed_reg[0]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[0]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[16]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[24]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[32]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[40]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[48]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[56]_i_1_n_9 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_0 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_1 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_10 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_11 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_12 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_13 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_14 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_15 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_2 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_3 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_4 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_5 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_6 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_7 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_8 ;
  wire \multicast_frame_transed_reg[8]_i_1_n_9 ;
  wire \multicast_received_good[0]_i_2_n_0 ;
  wire [63:0]multicast_received_good_reg;
  wire \multicast_received_good_reg[0]_i_1_n_0 ;
  wire \multicast_received_good_reg[0]_i_1_n_1 ;
  wire \multicast_received_good_reg[0]_i_1_n_10 ;
  wire \multicast_received_good_reg[0]_i_1_n_11 ;
  wire \multicast_received_good_reg[0]_i_1_n_12 ;
  wire \multicast_received_good_reg[0]_i_1_n_13 ;
  wire \multicast_received_good_reg[0]_i_1_n_14 ;
  wire \multicast_received_good_reg[0]_i_1_n_15 ;
  wire \multicast_received_good_reg[0]_i_1_n_2 ;
  wire \multicast_received_good_reg[0]_i_1_n_3 ;
  wire \multicast_received_good_reg[0]_i_1_n_4 ;
  wire \multicast_received_good_reg[0]_i_1_n_5 ;
  wire \multicast_received_good_reg[0]_i_1_n_6 ;
  wire \multicast_received_good_reg[0]_i_1_n_7 ;
  wire \multicast_received_good_reg[0]_i_1_n_8 ;
  wire \multicast_received_good_reg[0]_i_1_n_9 ;
  wire \multicast_received_good_reg[16]_i_1_n_0 ;
  wire \multicast_received_good_reg[16]_i_1_n_1 ;
  wire \multicast_received_good_reg[16]_i_1_n_10 ;
  wire \multicast_received_good_reg[16]_i_1_n_11 ;
  wire \multicast_received_good_reg[16]_i_1_n_12 ;
  wire \multicast_received_good_reg[16]_i_1_n_13 ;
  wire \multicast_received_good_reg[16]_i_1_n_14 ;
  wire \multicast_received_good_reg[16]_i_1_n_15 ;
  wire \multicast_received_good_reg[16]_i_1_n_2 ;
  wire \multicast_received_good_reg[16]_i_1_n_3 ;
  wire \multicast_received_good_reg[16]_i_1_n_4 ;
  wire \multicast_received_good_reg[16]_i_1_n_5 ;
  wire \multicast_received_good_reg[16]_i_1_n_6 ;
  wire \multicast_received_good_reg[16]_i_1_n_7 ;
  wire \multicast_received_good_reg[16]_i_1_n_8 ;
  wire \multicast_received_good_reg[16]_i_1_n_9 ;
  wire \multicast_received_good_reg[24]_i_1_n_0 ;
  wire \multicast_received_good_reg[24]_i_1_n_1 ;
  wire \multicast_received_good_reg[24]_i_1_n_10 ;
  wire \multicast_received_good_reg[24]_i_1_n_11 ;
  wire \multicast_received_good_reg[24]_i_1_n_12 ;
  wire \multicast_received_good_reg[24]_i_1_n_13 ;
  wire \multicast_received_good_reg[24]_i_1_n_14 ;
  wire \multicast_received_good_reg[24]_i_1_n_15 ;
  wire \multicast_received_good_reg[24]_i_1_n_2 ;
  wire \multicast_received_good_reg[24]_i_1_n_3 ;
  wire \multicast_received_good_reg[24]_i_1_n_4 ;
  wire \multicast_received_good_reg[24]_i_1_n_5 ;
  wire \multicast_received_good_reg[24]_i_1_n_6 ;
  wire \multicast_received_good_reg[24]_i_1_n_7 ;
  wire \multicast_received_good_reg[24]_i_1_n_8 ;
  wire \multicast_received_good_reg[24]_i_1_n_9 ;
  wire \multicast_received_good_reg[32]_i_1_n_0 ;
  wire \multicast_received_good_reg[32]_i_1_n_1 ;
  wire \multicast_received_good_reg[32]_i_1_n_10 ;
  wire \multicast_received_good_reg[32]_i_1_n_11 ;
  wire \multicast_received_good_reg[32]_i_1_n_12 ;
  wire \multicast_received_good_reg[32]_i_1_n_13 ;
  wire \multicast_received_good_reg[32]_i_1_n_14 ;
  wire \multicast_received_good_reg[32]_i_1_n_15 ;
  wire \multicast_received_good_reg[32]_i_1_n_2 ;
  wire \multicast_received_good_reg[32]_i_1_n_3 ;
  wire \multicast_received_good_reg[32]_i_1_n_4 ;
  wire \multicast_received_good_reg[32]_i_1_n_5 ;
  wire \multicast_received_good_reg[32]_i_1_n_6 ;
  wire \multicast_received_good_reg[32]_i_1_n_7 ;
  wire \multicast_received_good_reg[32]_i_1_n_8 ;
  wire \multicast_received_good_reg[32]_i_1_n_9 ;
  wire \multicast_received_good_reg[40]_i_1_n_0 ;
  wire \multicast_received_good_reg[40]_i_1_n_1 ;
  wire \multicast_received_good_reg[40]_i_1_n_10 ;
  wire \multicast_received_good_reg[40]_i_1_n_11 ;
  wire \multicast_received_good_reg[40]_i_1_n_12 ;
  wire \multicast_received_good_reg[40]_i_1_n_13 ;
  wire \multicast_received_good_reg[40]_i_1_n_14 ;
  wire \multicast_received_good_reg[40]_i_1_n_15 ;
  wire \multicast_received_good_reg[40]_i_1_n_2 ;
  wire \multicast_received_good_reg[40]_i_1_n_3 ;
  wire \multicast_received_good_reg[40]_i_1_n_4 ;
  wire \multicast_received_good_reg[40]_i_1_n_5 ;
  wire \multicast_received_good_reg[40]_i_1_n_6 ;
  wire \multicast_received_good_reg[40]_i_1_n_7 ;
  wire \multicast_received_good_reg[40]_i_1_n_8 ;
  wire \multicast_received_good_reg[40]_i_1_n_9 ;
  wire \multicast_received_good_reg[48]_i_1_n_0 ;
  wire \multicast_received_good_reg[48]_i_1_n_1 ;
  wire \multicast_received_good_reg[48]_i_1_n_10 ;
  wire \multicast_received_good_reg[48]_i_1_n_11 ;
  wire \multicast_received_good_reg[48]_i_1_n_12 ;
  wire \multicast_received_good_reg[48]_i_1_n_13 ;
  wire \multicast_received_good_reg[48]_i_1_n_14 ;
  wire \multicast_received_good_reg[48]_i_1_n_15 ;
  wire \multicast_received_good_reg[48]_i_1_n_2 ;
  wire \multicast_received_good_reg[48]_i_1_n_3 ;
  wire \multicast_received_good_reg[48]_i_1_n_4 ;
  wire \multicast_received_good_reg[48]_i_1_n_5 ;
  wire \multicast_received_good_reg[48]_i_1_n_6 ;
  wire \multicast_received_good_reg[48]_i_1_n_7 ;
  wire \multicast_received_good_reg[48]_i_1_n_8 ;
  wire \multicast_received_good_reg[48]_i_1_n_9 ;
  wire \multicast_received_good_reg[56]_i_1_n_1 ;
  wire \multicast_received_good_reg[56]_i_1_n_10 ;
  wire \multicast_received_good_reg[56]_i_1_n_11 ;
  wire \multicast_received_good_reg[56]_i_1_n_12 ;
  wire \multicast_received_good_reg[56]_i_1_n_13 ;
  wire \multicast_received_good_reg[56]_i_1_n_14 ;
  wire \multicast_received_good_reg[56]_i_1_n_15 ;
  wire \multicast_received_good_reg[56]_i_1_n_2 ;
  wire \multicast_received_good_reg[56]_i_1_n_3 ;
  wire \multicast_received_good_reg[56]_i_1_n_4 ;
  wire \multicast_received_good_reg[56]_i_1_n_5 ;
  wire \multicast_received_good_reg[56]_i_1_n_6 ;
  wire \multicast_received_good_reg[56]_i_1_n_7 ;
  wire \multicast_received_good_reg[56]_i_1_n_8 ;
  wire \multicast_received_good_reg[56]_i_1_n_9 ;
  wire \multicast_received_good_reg[8]_i_1_n_0 ;
  wire \multicast_received_good_reg[8]_i_1_n_1 ;
  wire \multicast_received_good_reg[8]_i_1_n_10 ;
  wire \multicast_received_good_reg[8]_i_1_n_11 ;
  wire \multicast_received_good_reg[8]_i_1_n_12 ;
  wire \multicast_received_good_reg[8]_i_1_n_13 ;
  wire \multicast_received_good_reg[8]_i_1_n_14 ;
  wire \multicast_received_good_reg[8]_i_1_n_15 ;
  wire \multicast_received_good_reg[8]_i_1_n_2 ;
  wire \multicast_received_good_reg[8]_i_1_n_3 ;
  wire \multicast_received_good_reg[8]_i_1_n_4 ;
  wire \multicast_received_good_reg[8]_i_1_n_5 ;
  wire \multicast_received_good_reg[8]_i_1_n_6 ;
  wire \multicast_received_good_reg[8]_i_1_n_7 ;
  wire \multicast_received_good_reg[8]_i_1_n_8 ;
  wire \multicast_received_good_reg[8]_i_1_n_9 ;
  wire [9:0]out;
  wire \oversize_frame_good[0]_i_2_n_0 ;
  wire [63:0]oversize_frame_good_reg;
  wire \oversize_frame_good_reg[0]_i_1_n_0 ;
  wire \oversize_frame_good_reg[0]_i_1_n_1 ;
  wire \oversize_frame_good_reg[0]_i_1_n_10 ;
  wire \oversize_frame_good_reg[0]_i_1_n_11 ;
  wire \oversize_frame_good_reg[0]_i_1_n_12 ;
  wire \oversize_frame_good_reg[0]_i_1_n_13 ;
  wire \oversize_frame_good_reg[0]_i_1_n_14 ;
  wire \oversize_frame_good_reg[0]_i_1_n_15 ;
  wire \oversize_frame_good_reg[0]_i_1_n_2 ;
  wire \oversize_frame_good_reg[0]_i_1_n_3 ;
  wire \oversize_frame_good_reg[0]_i_1_n_4 ;
  wire \oversize_frame_good_reg[0]_i_1_n_5 ;
  wire \oversize_frame_good_reg[0]_i_1_n_6 ;
  wire \oversize_frame_good_reg[0]_i_1_n_7 ;
  wire \oversize_frame_good_reg[0]_i_1_n_8 ;
  wire \oversize_frame_good_reg[0]_i_1_n_9 ;
  wire \oversize_frame_good_reg[16]_i_1_n_0 ;
  wire \oversize_frame_good_reg[16]_i_1_n_1 ;
  wire \oversize_frame_good_reg[16]_i_1_n_10 ;
  wire \oversize_frame_good_reg[16]_i_1_n_11 ;
  wire \oversize_frame_good_reg[16]_i_1_n_12 ;
  wire \oversize_frame_good_reg[16]_i_1_n_13 ;
  wire \oversize_frame_good_reg[16]_i_1_n_14 ;
  wire \oversize_frame_good_reg[16]_i_1_n_15 ;
  wire \oversize_frame_good_reg[16]_i_1_n_2 ;
  wire \oversize_frame_good_reg[16]_i_1_n_3 ;
  wire \oversize_frame_good_reg[16]_i_1_n_4 ;
  wire \oversize_frame_good_reg[16]_i_1_n_5 ;
  wire \oversize_frame_good_reg[16]_i_1_n_6 ;
  wire \oversize_frame_good_reg[16]_i_1_n_7 ;
  wire \oversize_frame_good_reg[16]_i_1_n_8 ;
  wire \oversize_frame_good_reg[16]_i_1_n_9 ;
  wire \oversize_frame_good_reg[24]_i_1_n_0 ;
  wire \oversize_frame_good_reg[24]_i_1_n_1 ;
  wire \oversize_frame_good_reg[24]_i_1_n_10 ;
  wire \oversize_frame_good_reg[24]_i_1_n_11 ;
  wire \oversize_frame_good_reg[24]_i_1_n_12 ;
  wire \oversize_frame_good_reg[24]_i_1_n_13 ;
  wire \oversize_frame_good_reg[24]_i_1_n_14 ;
  wire \oversize_frame_good_reg[24]_i_1_n_15 ;
  wire \oversize_frame_good_reg[24]_i_1_n_2 ;
  wire \oversize_frame_good_reg[24]_i_1_n_3 ;
  wire \oversize_frame_good_reg[24]_i_1_n_4 ;
  wire \oversize_frame_good_reg[24]_i_1_n_5 ;
  wire \oversize_frame_good_reg[24]_i_1_n_6 ;
  wire \oversize_frame_good_reg[24]_i_1_n_7 ;
  wire \oversize_frame_good_reg[24]_i_1_n_8 ;
  wire \oversize_frame_good_reg[24]_i_1_n_9 ;
  wire \oversize_frame_good_reg[32]_i_1_n_0 ;
  wire \oversize_frame_good_reg[32]_i_1_n_1 ;
  wire \oversize_frame_good_reg[32]_i_1_n_10 ;
  wire \oversize_frame_good_reg[32]_i_1_n_11 ;
  wire \oversize_frame_good_reg[32]_i_1_n_12 ;
  wire \oversize_frame_good_reg[32]_i_1_n_13 ;
  wire \oversize_frame_good_reg[32]_i_1_n_14 ;
  wire \oversize_frame_good_reg[32]_i_1_n_15 ;
  wire \oversize_frame_good_reg[32]_i_1_n_2 ;
  wire \oversize_frame_good_reg[32]_i_1_n_3 ;
  wire \oversize_frame_good_reg[32]_i_1_n_4 ;
  wire \oversize_frame_good_reg[32]_i_1_n_5 ;
  wire \oversize_frame_good_reg[32]_i_1_n_6 ;
  wire \oversize_frame_good_reg[32]_i_1_n_7 ;
  wire \oversize_frame_good_reg[32]_i_1_n_8 ;
  wire \oversize_frame_good_reg[32]_i_1_n_9 ;
  wire \oversize_frame_good_reg[40]_i_1_n_0 ;
  wire \oversize_frame_good_reg[40]_i_1_n_1 ;
  wire \oversize_frame_good_reg[40]_i_1_n_10 ;
  wire \oversize_frame_good_reg[40]_i_1_n_11 ;
  wire \oversize_frame_good_reg[40]_i_1_n_12 ;
  wire \oversize_frame_good_reg[40]_i_1_n_13 ;
  wire \oversize_frame_good_reg[40]_i_1_n_14 ;
  wire \oversize_frame_good_reg[40]_i_1_n_15 ;
  wire \oversize_frame_good_reg[40]_i_1_n_2 ;
  wire \oversize_frame_good_reg[40]_i_1_n_3 ;
  wire \oversize_frame_good_reg[40]_i_1_n_4 ;
  wire \oversize_frame_good_reg[40]_i_1_n_5 ;
  wire \oversize_frame_good_reg[40]_i_1_n_6 ;
  wire \oversize_frame_good_reg[40]_i_1_n_7 ;
  wire \oversize_frame_good_reg[40]_i_1_n_8 ;
  wire \oversize_frame_good_reg[40]_i_1_n_9 ;
  wire \oversize_frame_good_reg[48]_i_1_n_0 ;
  wire \oversize_frame_good_reg[48]_i_1_n_1 ;
  wire \oversize_frame_good_reg[48]_i_1_n_10 ;
  wire \oversize_frame_good_reg[48]_i_1_n_11 ;
  wire \oversize_frame_good_reg[48]_i_1_n_12 ;
  wire \oversize_frame_good_reg[48]_i_1_n_13 ;
  wire \oversize_frame_good_reg[48]_i_1_n_14 ;
  wire \oversize_frame_good_reg[48]_i_1_n_15 ;
  wire \oversize_frame_good_reg[48]_i_1_n_2 ;
  wire \oversize_frame_good_reg[48]_i_1_n_3 ;
  wire \oversize_frame_good_reg[48]_i_1_n_4 ;
  wire \oversize_frame_good_reg[48]_i_1_n_5 ;
  wire \oversize_frame_good_reg[48]_i_1_n_6 ;
  wire \oversize_frame_good_reg[48]_i_1_n_7 ;
  wire \oversize_frame_good_reg[48]_i_1_n_8 ;
  wire \oversize_frame_good_reg[48]_i_1_n_9 ;
  wire \oversize_frame_good_reg[56]_i_1_n_1 ;
  wire \oversize_frame_good_reg[56]_i_1_n_10 ;
  wire \oversize_frame_good_reg[56]_i_1_n_11 ;
  wire \oversize_frame_good_reg[56]_i_1_n_12 ;
  wire \oversize_frame_good_reg[56]_i_1_n_13 ;
  wire \oversize_frame_good_reg[56]_i_1_n_14 ;
  wire \oversize_frame_good_reg[56]_i_1_n_15 ;
  wire \oversize_frame_good_reg[56]_i_1_n_2 ;
  wire \oversize_frame_good_reg[56]_i_1_n_3 ;
  wire \oversize_frame_good_reg[56]_i_1_n_4 ;
  wire \oversize_frame_good_reg[56]_i_1_n_5 ;
  wire \oversize_frame_good_reg[56]_i_1_n_6 ;
  wire \oversize_frame_good_reg[56]_i_1_n_7 ;
  wire \oversize_frame_good_reg[56]_i_1_n_8 ;
  wire \oversize_frame_good_reg[56]_i_1_n_9 ;
  wire \oversize_frame_good_reg[8]_i_1_n_0 ;
  wire \oversize_frame_good_reg[8]_i_1_n_1 ;
  wire \oversize_frame_good_reg[8]_i_1_n_10 ;
  wire \oversize_frame_good_reg[8]_i_1_n_11 ;
  wire \oversize_frame_good_reg[8]_i_1_n_12 ;
  wire \oversize_frame_good_reg[8]_i_1_n_13 ;
  wire \oversize_frame_good_reg[8]_i_1_n_14 ;
  wire \oversize_frame_good_reg[8]_i_1_n_15 ;
  wire \oversize_frame_good_reg[8]_i_1_n_2 ;
  wire \oversize_frame_good_reg[8]_i_1_n_3 ;
  wire \oversize_frame_good_reg[8]_i_1_n_4 ;
  wire \oversize_frame_good_reg[8]_i_1_n_5 ;
  wire \oversize_frame_good_reg[8]_i_1_n_6 ;
  wire \oversize_frame_good_reg[8]_i_1_n_7 ;
  wire \oversize_frame_good_reg[8]_i_1_n_8 ;
  wire \oversize_frame_good_reg[8]_i_1_n_9 ;
  wire \oversize_frame_transed[0]_i_2_n_0 ;
  wire [63:0]oversize_frame_transed_reg;
  wire \oversize_frame_transed_reg[0]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[0]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[16]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[24]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[32]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[40]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[48]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[56]_i_1_n_9 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_0 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_1 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_10 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_11 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_12 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_13 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_14 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_15 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_2 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_3 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_4 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_5 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_6 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_7 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_8 ;
  wire \oversize_frame_transed_reg[8]_i_1_n_9 ;
  wire [63:0]p_0_in;
  wire [31:0]p_1_in;
  wire \pause_frame_good[0]_i_2_n_0 ;
  wire [63:0]pause_frame_good_reg;
  wire \pause_frame_good_reg[0]_i_1_n_0 ;
  wire \pause_frame_good_reg[0]_i_1_n_1 ;
  wire \pause_frame_good_reg[0]_i_1_n_10 ;
  wire \pause_frame_good_reg[0]_i_1_n_11 ;
  wire \pause_frame_good_reg[0]_i_1_n_12 ;
  wire \pause_frame_good_reg[0]_i_1_n_13 ;
  wire \pause_frame_good_reg[0]_i_1_n_14 ;
  wire \pause_frame_good_reg[0]_i_1_n_15 ;
  wire \pause_frame_good_reg[0]_i_1_n_2 ;
  wire \pause_frame_good_reg[0]_i_1_n_3 ;
  wire \pause_frame_good_reg[0]_i_1_n_4 ;
  wire \pause_frame_good_reg[0]_i_1_n_5 ;
  wire \pause_frame_good_reg[0]_i_1_n_6 ;
  wire \pause_frame_good_reg[0]_i_1_n_7 ;
  wire \pause_frame_good_reg[0]_i_1_n_8 ;
  wire \pause_frame_good_reg[0]_i_1_n_9 ;
  wire \pause_frame_good_reg[16]_i_1_n_0 ;
  wire \pause_frame_good_reg[16]_i_1_n_1 ;
  wire \pause_frame_good_reg[16]_i_1_n_10 ;
  wire \pause_frame_good_reg[16]_i_1_n_11 ;
  wire \pause_frame_good_reg[16]_i_1_n_12 ;
  wire \pause_frame_good_reg[16]_i_1_n_13 ;
  wire \pause_frame_good_reg[16]_i_1_n_14 ;
  wire \pause_frame_good_reg[16]_i_1_n_15 ;
  wire \pause_frame_good_reg[16]_i_1_n_2 ;
  wire \pause_frame_good_reg[16]_i_1_n_3 ;
  wire \pause_frame_good_reg[16]_i_1_n_4 ;
  wire \pause_frame_good_reg[16]_i_1_n_5 ;
  wire \pause_frame_good_reg[16]_i_1_n_6 ;
  wire \pause_frame_good_reg[16]_i_1_n_7 ;
  wire \pause_frame_good_reg[16]_i_1_n_8 ;
  wire \pause_frame_good_reg[16]_i_1_n_9 ;
  wire \pause_frame_good_reg[24]_i_1_n_0 ;
  wire \pause_frame_good_reg[24]_i_1_n_1 ;
  wire \pause_frame_good_reg[24]_i_1_n_10 ;
  wire \pause_frame_good_reg[24]_i_1_n_11 ;
  wire \pause_frame_good_reg[24]_i_1_n_12 ;
  wire \pause_frame_good_reg[24]_i_1_n_13 ;
  wire \pause_frame_good_reg[24]_i_1_n_14 ;
  wire \pause_frame_good_reg[24]_i_1_n_15 ;
  wire \pause_frame_good_reg[24]_i_1_n_2 ;
  wire \pause_frame_good_reg[24]_i_1_n_3 ;
  wire \pause_frame_good_reg[24]_i_1_n_4 ;
  wire \pause_frame_good_reg[24]_i_1_n_5 ;
  wire \pause_frame_good_reg[24]_i_1_n_6 ;
  wire \pause_frame_good_reg[24]_i_1_n_7 ;
  wire \pause_frame_good_reg[24]_i_1_n_8 ;
  wire \pause_frame_good_reg[24]_i_1_n_9 ;
  wire \pause_frame_good_reg[32]_i_1_n_0 ;
  wire \pause_frame_good_reg[32]_i_1_n_1 ;
  wire \pause_frame_good_reg[32]_i_1_n_10 ;
  wire \pause_frame_good_reg[32]_i_1_n_11 ;
  wire \pause_frame_good_reg[32]_i_1_n_12 ;
  wire \pause_frame_good_reg[32]_i_1_n_13 ;
  wire \pause_frame_good_reg[32]_i_1_n_14 ;
  wire \pause_frame_good_reg[32]_i_1_n_15 ;
  wire \pause_frame_good_reg[32]_i_1_n_2 ;
  wire \pause_frame_good_reg[32]_i_1_n_3 ;
  wire \pause_frame_good_reg[32]_i_1_n_4 ;
  wire \pause_frame_good_reg[32]_i_1_n_5 ;
  wire \pause_frame_good_reg[32]_i_1_n_6 ;
  wire \pause_frame_good_reg[32]_i_1_n_7 ;
  wire \pause_frame_good_reg[32]_i_1_n_8 ;
  wire \pause_frame_good_reg[32]_i_1_n_9 ;
  wire \pause_frame_good_reg[40]_i_1_n_0 ;
  wire \pause_frame_good_reg[40]_i_1_n_1 ;
  wire \pause_frame_good_reg[40]_i_1_n_10 ;
  wire \pause_frame_good_reg[40]_i_1_n_11 ;
  wire \pause_frame_good_reg[40]_i_1_n_12 ;
  wire \pause_frame_good_reg[40]_i_1_n_13 ;
  wire \pause_frame_good_reg[40]_i_1_n_14 ;
  wire \pause_frame_good_reg[40]_i_1_n_15 ;
  wire \pause_frame_good_reg[40]_i_1_n_2 ;
  wire \pause_frame_good_reg[40]_i_1_n_3 ;
  wire \pause_frame_good_reg[40]_i_1_n_4 ;
  wire \pause_frame_good_reg[40]_i_1_n_5 ;
  wire \pause_frame_good_reg[40]_i_1_n_6 ;
  wire \pause_frame_good_reg[40]_i_1_n_7 ;
  wire \pause_frame_good_reg[40]_i_1_n_8 ;
  wire \pause_frame_good_reg[40]_i_1_n_9 ;
  wire \pause_frame_good_reg[48]_i_1_n_0 ;
  wire \pause_frame_good_reg[48]_i_1_n_1 ;
  wire \pause_frame_good_reg[48]_i_1_n_10 ;
  wire \pause_frame_good_reg[48]_i_1_n_11 ;
  wire \pause_frame_good_reg[48]_i_1_n_12 ;
  wire \pause_frame_good_reg[48]_i_1_n_13 ;
  wire \pause_frame_good_reg[48]_i_1_n_14 ;
  wire \pause_frame_good_reg[48]_i_1_n_15 ;
  wire \pause_frame_good_reg[48]_i_1_n_2 ;
  wire \pause_frame_good_reg[48]_i_1_n_3 ;
  wire \pause_frame_good_reg[48]_i_1_n_4 ;
  wire \pause_frame_good_reg[48]_i_1_n_5 ;
  wire \pause_frame_good_reg[48]_i_1_n_6 ;
  wire \pause_frame_good_reg[48]_i_1_n_7 ;
  wire \pause_frame_good_reg[48]_i_1_n_8 ;
  wire \pause_frame_good_reg[48]_i_1_n_9 ;
  wire \pause_frame_good_reg[56]_i_1_n_1 ;
  wire \pause_frame_good_reg[56]_i_1_n_10 ;
  wire \pause_frame_good_reg[56]_i_1_n_11 ;
  wire \pause_frame_good_reg[56]_i_1_n_12 ;
  wire \pause_frame_good_reg[56]_i_1_n_13 ;
  wire \pause_frame_good_reg[56]_i_1_n_14 ;
  wire \pause_frame_good_reg[56]_i_1_n_15 ;
  wire \pause_frame_good_reg[56]_i_1_n_2 ;
  wire \pause_frame_good_reg[56]_i_1_n_3 ;
  wire \pause_frame_good_reg[56]_i_1_n_4 ;
  wire \pause_frame_good_reg[56]_i_1_n_5 ;
  wire \pause_frame_good_reg[56]_i_1_n_6 ;
  wire \pause_frame_good_reg[56]_i_1_n_7 ;
  wire \pause_frame_good_reg[56]_i_1_n_8 ;
  wire \pause_frame_good_reg[56]_i_1_n_9 ;
  wire \pause_frame_good_reg[8]_i_1_n_0 ;
  wire \pause_frame_good_reg[8]_i_1_n_1 ;
  wire \pause_frame_good_reg[8]_i_1_n_10 ;
  wire \pause_frame_good_reg[8]_i_1_n_11 ;
  wire \pause_frame_good_reg[8]_i_1_n_12 ;
  wire \pause_frame_good_reg[8]_i_1_n_13 ;
  wire \pause_frame_good_reg[8]_i_1_n_14 ;
  wire \pause_frame_good_reg[8]_i_1_n_15 ;
  wire \pause_frame_good_reg[8]_i_1_n_2 ;
  wire \pause_frame_good_reg[8]_i_1_n_3 ;
  wire \pause_frame_good_reg[8]_i_1_n_4 ;
  wire \pause_frame_good_reg[8]_i_1_n_5 ;
  wire \pause_frame_good_reg[8]_i_1_n_6 ;
  wire \pause_frame_good_reg[8]_i_1_n_7 ;
  wire \pause_frame_good_reg[8]_i_1_n_8 ;
  wire \pause_frame_good_reg[8]_i_1_n_9 ;
  wire \pause_frame_transed[0]_i_2_n_0 ;
  wire [63:0]pause_frame_transed_reg;
  wire \pause_frame_transed_reg[0]_i_1_n_0 ;
  wire \pause_frame_transed_reg[0]_i_1_n_1 ;
  wire \pause_frame_transed_reg[0]_i_1_n_10 ;
  wire \pause_frame_transed_reg[0]_i_1_n_11 ;
  wire \pause_frame_transed_reg[0]_i_1_n_12 ;
  wire \pause_frame_transed_reg[0]_i_1_n_13 ;
  wire \pause_frame_transed_reg[0]_i_1_n_14 ;
  wire \pause_frame_transed_reg[0]_i_1_n_15 ;
  wire \pause_frame_transed_reg[0]_i_1_n_2 ;
  wire \pause_frame_transed_reg[0]_i_1_n_3 ;
  wire \pause_frame_transed_reg[0]_i_1_n_4 ;
  wire \pause_frame_transed_reg[0]_i_1_n_5 ;
  wire \pause_frame_transed_reg[0]_i_1_n_6 ;
  wire \pause_frame_transed_reg[0]_i_1_n_7 ;
  wire \pause_frame_transed_reg[0]_i_1_n_8 ;
  wire \pause_frame_transed_reg[0]_i_1_n_9 ;
  wire \pause_frame_transed_reg[16]_i_1_n_0 ;
  wire \pause_frame_transed_reg[16]_i_1_n_1 ;
  wire \pause_frame_transed_reg[16]_i_1_n_10 ;
  wire \pause_frame_transed_reg[16]_i_1_n_11 ;
  wire \pause_frame_transed_reg[16]_i_1_n_12 ;
  wire \pause_frame_transed_reg[16]_i_1_n_13 ;
  wire \pause_frame_transed_reg[16]_i_1_n_14 ;
  wire \pause_frame_transed_reg[16]_i_1_n_15 ;
  wire \pause_frame_transed_reg[16]_i_1_n_2 ;
  wire \pause_frame_transed_reg[16]_i_1_n_3 ;
  wire \pause_frame_transed_reg[16]_i_1_n_4 ;
  wire \pause_frame_transed_reg[16]_i_1_n_5 ;
  wire \pause_frame_transed_reg[16]_i_1_n_6 ;
  wire \pause_frame_transed_reg[16]_i_1_n_7 ;
  wire \pause_frame_transed_reg[16]_i_1_n_8 ;
  wire \pause_frame_transed_reg[16]_i_1_n_9 ;
  wire \pause_frame_transed_reg[24]_i_1_n_0 ;
  wire \pause_frame_transed_reg[24]_i_1_n_1 ;
  wire \pause_frame_transed_reg[24]_i_1_n_10 ;
  wire \pause_frame_transed_reg[24]_i_1_n_11 ;
  wire \pause_frame_transed_reg[24]_i_1_n_12 ;
  wire \pause_frame_transed_reg[24]_i_1_n_13 ;
  wire \pause_frame_transed_reg[24]_i_1_n_14 ;
  wire \pause_frame_transed_reg[24]_i_1_n_15 ;
  wire \pause_frame_transed_reg[24]_i_1_n_2 ;
  wire \pause_frame_transed_reg[24]_i_1_n_3 ;
  wire \pause_frame_transed_reg[24]_i_1_n_4 ;
  wire \pause_frame_transed_reg[24]_i_1_n_5 ;
  wire \pause_frame_transed_reg[24]_i_1_n_6 ;
  wire \pause_frame_transed_reg[24]_i_1_n_7 ;
  wire \pause_frame_transed_reg[24]_i_1_n_8 ;
  wire \pause_frame_transed_reg[24]_i_1_n_9 ;
  wire \pause_frame_transed_reg[32]_i_1_n_0 ;
  wire \pause_frame_transed_reg[32]_i_1_n_1 ;
  wire \pause_frame_transed_reg[32]_i_1_n_10 ;
  wire \pause_frame_transed_reg[32]_i_1_n_11 ;
  wire \pause_frame_transed_reg[32]_i_1_n_12 ;
  wire \pause_frame_transed_reg[32]_i_1_n_13 ;
  wire \pause_frame_transed_reg[32]_i_1_n_14 ;
  wire \pause_frame_transed_reg[32]_i_1_n_15 ;
  wire \pause_frame_transed_reg[32]_i_1_n_2 ;
  wire \pause_frame_transed_reg[32]_i_1_n_3 ;
  wire \pause_frame_transed_reg[32]_i_1_n_4 ;
  wire \pause_frame_transed_reg[32]_i_1_n_5 ;
  wire \pause_frame_transed_reg[32]_i_1_n_6 ;
  wire \pause_frame_transed_reg[32]_i_1_n_7 ;
  wire \pause_frame_transed_reg[32]_i_1_n_8 ;
  wire \pause_frame_transed_reg[32]_i_1_n_9 ;
  wire \pause_frame_transed_reg[40]_i_1_n_0 ;
  wire \pause_frame_transed_reg[40]_i_1_n_1 ;
  wire \pause_frame_transed_reg[40]_i_1_n_10 ;
  wire \pause_frame_transed_reg[40]_i_1_n_11 ;
  wire \pause_frame_transed_reg[40]_i_1_n_12 ;
  wire \pause_frame_transed_reg[40]_i_1_n_13 ;
  wire \pause_frame_transed_reg[40]_i_1_n_14 ;
  wire \pause_frame_transed_reg[40]_i_1_n_15 ;
  wire \pause_frame_transed_reg[40]_i_1_n_2 ;
  wire \pause_frame_transed_reg[40]_i_1_n_3 ;
  wire \pause_frame_transed_reg[40]_i_1_n_4 ;
  wire \pause_frame_transed_reg[40]_i_1_n_5 ;
  wire \pause_frame_transed_reg[40]_i_1_n_6 ;
  wire \pause_frame_transed_reg[40]_i_1_n_7 ;
  wire \pause_frame_transed_reg[40]_i_1_n_8 ;
  wire \pause_frame_transed_reg[40]_i_1_n_9 ;
  wire \pause_frame_transed_reg[48]_i_1_n_0 ;
  wire \pause_frame_transed_reg[48]_i_1_n_1 ;
  wire \pause_frame_transed_reg[48]_i_1_n_10 ;
  wire \pause_frame_transed_reg[48]_i_1_n_11 ;
  wire \pause_frame_transed_reg[48]_i_1_n_12 ;
  wire \pause_frame_transed_reg[48]_i_1_n_13 ;
  wire \pause_frame_transed_reg[48]_i_1_n_14 ;
  wire \pause_frame_transed_reg[48]_i_1_n_15 ;
  wire \pause_frame_transed_reg[48]_i_1_n_2 ;
  wire \pause_frame_transed_reg[48]_i_1_n_3 ;
  wire \pause_frame_transed_reg[48]_i_1_n_4 ;
  wire \pause_frame_transed_reg[48]_i_1_n_5 ;
  wire \pause_frame_transed_reg[48]_i_1_n_6 ;
  wire \pause_frame_transed_reg[48]_i_1_n_7 ;
  wire \pause_frame_transed_reg[48]_i_1_n_8 ;
  wire \pause_frame_transed_reg[48]_i_1_n_9 ;
  wire \pause_frame_transed_reg[56]_i_1_n_1 ;
  wire \pause_frame_transed_reg[56]_i_1_n_10 ;
  wire \pause_frame_transed_reg[56]_i_1_n_11 ;
  wire \pause_frame_transed_reg[56]_i_1_n_12 ;
  wire \pause_frame_transed_reg[56]_i_1_n_13 ;
  wire \pause_frame_transed_reg[56]_i_1_n_14 ;
  wire \pause_frame_transed_reg[56]_i_1_n_15 ;
  wire \pause_frame_transed_reg[56]_i_1_n_2 ;
  wire \pause_frame_transed_reg[56]_i_1_n_3 ;
  wire \pause_frame_transed_reg[56]_i_1_n_4 ;
  wire \pause_frame_transed_reg[56]_i_1_n_5 ;
  wire \pause_frame_transed_reg[56]_i_1_n_6 ;
  wire \pause_frame_transed_reg[56]_i_1_n_7 ;
  wire \pause_frame_transed_reg[56]_i_1_n_8 ;
  wire \pause_frame_transed_reg[56]_i_1_n_9 ;
  wire \pause_frame_transed_reg[8]_i_1_n_0 ;
  wire \pause_frame_transed_reg[8]_i_1_n_1 ;
  wire \pause_frame_transed_reg[8]_i_1_n_10 ;
  wire \pause_frame_transed_reg[8]_i_1_n_11 ;
  wire \pause_frame_transed_reg[8]_i_1_n_12 ;
  wire \pause_frame_transed_reg[8]_i_1_n_13 ;
  wire \pause_frame_transed_reg[8]_i_1_n_14 ;
  wire \pause_frame_transed_reg[8]_i_1_n_15 ;
  wire \pause_frame_transed_reg[8]_i_1_n_2 ;
  wire \pause_frame_transed_reg[8]_i_1_n_3 ;
  wire \pause_frame_transed_reg[8]_i_1_n_4 ;
  wire \pause_frame_transed_reg[8]_i_1_n_5 ;
  wire \pause_frame_transed_reg[8]_i_1_n_6 ;
  wire \pause_frame_transed_reg[8]_i_1_n_7 ;
  wire \pause_frame_transed_reg[8]_i_1_n_8 ;
  wire \pause_frame_transed_reg[8]_i_1_n_9 ;
  wire read_done;
  wire read_done_i_1_n_0;
  wire read_done_reg_n_0;
  wire recv_config01__0;
  wire \recv_config0[31]_i_1_n_0 ;
  wire \recv_config0[31]_i_2_n_0 ;
  wire \recv_config0[31]_i_3_n_0 ;
  wire [0:0]\recv_config0_reg[0]_0 ;
  wire \recv_config1[31]_i_1_n_0 ;
  wire \recv_config1[31]_i_3_n_0 ;
  wire \recv_config1[31]_i_4_n_0 ;
  wire \recv_config1_reg_n_0_[16] ;
  wire \recv_config1_reg_n_0_[17] ;
  wire \recv_config1_reg_n_0_[18] ;
  wire \recv_config1_reg_n_0_[19] ;
  wire \recv_config1_reg_n_0_[20] ;
  wire \recv_config1_reg_n_0_[21] ;
  wire \recv_config1_reg_n_0_[22] ;
  wire \recv_config1_reg_n_0_[23] ;
  wire \recv_config1_reg_n_0_[24] ;
  wire \recv_config1_reg_n_0_[25] ;
  wire \recv_config1_reg_n_0_[26] ;
  wire \rs_config[31]_i_1_n_0 ;
  wire \rs_config[31]_i_2_n_0 ;
  wire \rs_config_reg_n_0_[0] ;
  wire \rs_config_reg_n_0_[10] ;
  wire \rs_config_reg_n_0_[11] ;
  wire \rs_config_reg_n_0_[12] ;
  wire \rs_config_reg_n_0_[13] ;
  wire \rs_config_reg_n_0_[14] ;
  wire \rs_config_reg_n_0_[15] ;
  wire \rs_config_reg_n_0_[16] ;
  wire \rs_config_reg_n_0_[17] ;
  wire \rs_config_reg_n_0_[18] ;
  wire \rs_config_reg_n_0_[19] ;
  wire \rs_config_reg_n_0_[1] ;
  wire \rs_config_reg_n_0_[20] ;
  wire \rs_config_reg_n_0_[21] ;
  wire \rs_config_reg_n_0_[22] ;
  wire \rs_config_reg_n_0_[23] ;
  wire \rs_config_reg_n_0_[24] ;
  wire \rs_config_reg_n_0_[25] ;
  wire \rs_config_reg_n_0_[26] ;
  wire \rs_config_reg_n_0_[28] ;
  wire \rs_config_reg_n_0_[29] ;
  wire \rs_config_reg_n_0_[2] ;
  wire \rs_config_reg_n_0_[30] ;
  wire \rs_config_reg_n_0_[31] ;
  wire \rs_config_reg_n_0_[3] ;
  wire \rs_config_reg_n_0_[4] ;
  wire \rs_config_reg_n_0_[5] ;
  wire \rs_config_reg_n_0_[6] ;
  wire \rs_config_reg_n_0_[7] ;
  wire \rs_config_reg_n_0_[8] ;
  wire \rs_config_reg_n_0_[9] ;
  wire rst_i;
  wire [18:0]rxStatRegPlus;
  wire [4:0]sel0;
  wire [63:0]stat_rd_data;
  wire \stat_rd_data[0]_i_10_n_0 ;
  wire \stat_rd_data[0]_i_11_n_0 ;
  wire \stat_rd_data[0]_i_12_n_0 ;
  wire \stat_rd_data[0]_i_13_n_0 ;
  wire \stat_rd_data[0]_i_14_n_0 ;
  wire \stat_rd_data[0]_i_2_n_0 ;
  wire \stat_rd_data[0]_i_3_n_0 ;
  wire \stat_rd_data[0]_i_5_n_0 ;
  wire \stat_rd_data[0]_i_6_n_0 ;
  wire \stat_rd_data[0]_i_7_n_0 ;
  wire \stat_rd_data[10]_i_10_n_0 ;
  wire \stat_rd_data[10]_i_11_n_0 ;
  wire \stat_rd_data[10]_i_12_n_0 ;
  wire \stat_rd_data[10]_i_13_n_0 ;
  wire \stat_rd_data[10]_i_14_n_0 ;
  wire \stat_rd_data[10]_i_2_n_0 ;
  wire \stat_rd_data[10]_i_3_n_0 ;
  wire \stat_rd_data[10]_i_5_n_0 ;
  wire \stat_rd_data[10]_i_6_n_0 ;
  wire \stat_rd_data[10]_i_7_n_0 ;
  wire \stat_rd_data[11]_i_10_n_0 ;
  wire \stat_rd_data[11]_i_11_n_0 ;
  wire \stat_rd_data[11]_i_12_n_0 ;
  wire \stat_rd_data[11]_i_13_n_0 ;
  wire \stat_rd_data[11]_i_14_n_0 ;
  wire \stat_rd_data[11]_i_2_n_0 ;
  wire \stat_rd_data[11]_i_3_n_0 ;
  wire \stat_rd_data[11]_i_5_n_0 ;
  wire \stat_rd_data[11]_i_6_n_0 ;
  wire \stat_rd_data[11]_i_7_n_0 ;
  wire \stat_rd_data[12]_i_10_n_0 ;
  wire \stat_rd_data[12]_i_11_n_0 ;
  wire \stat_rd_data[12]_i_12_n_0 ;
  wire \stat_rd_data[12]_i_13_n_0 ;
  wire \stat_rd_data[12]_i_14_n_0 ;
  wire \stat_rd_data[12]_i_2_n_0 ;
  wire \stat_rd_data[12]_i_3_n_0 ;
  wire \stat_rd_data[12]_i_5_n_0 ;
  wire \stat_rd_data[12]_i_6_n_0 ;
  wire \stat_rd_data[12]_i_7_n_0 ;
  wire \stat_rd_data[13]_i_10_n_0 ;
  wire \stat_rd_data[13]_i_11_n_0 ;
  wire \stat_rd_data[13]_i_12_n_0 ;
  wire \stat_rd_data[13]_i_13_n_0 ;
  wire \stat_rd_data[13]_i_14_n_0 ;
  wire \stat_rd_data[13]_i_2_n_0 ;
  wire \stat_rd_data[13]_i_3_n_0 ;
  wire \stat_rd_data[13]_i_5_n_0 ;
  wire \stat_rd_data[13]_i_6_n_0 ;
  wire \stat_rd_data[13]_i_7_n_0 ;
  wire \stat_rd_data[14]_i_10_n_0 ;
  wire \stat_rd_data[14]_i_11_n_0 ;
  wire \stat_rd_data[14]_i_12_n_0 ;
  wire \stat_rd_data[14]_i_13_n_0 ;
  wire \stat_rd_data[14]_i_14_n_0 ;
  wire \stat_rd_data[14]_i_2_n_0 ;
  wire \stat_rd_data[14]_i_3_n_0 ;
  wire \stat_rd_data[14]_i_5_n_0 ;
  wire \stat_rd_data[14]_i_6_n_0 ;
  wire \stat_rd_data[14]_i_7_n_0 ;
  wire \stat_rd_data[15]_i_10_n_0 ;
  wire \stat_rd_data[15]_i_11_n_0 ;
  wire \stat_rd_data[15]_i_12_n_0 ;
  wire \stat_rd_data[15]_i_13_n_0 ;
  wire \stat_rd_data[15]_i_14_n_0 ;
  wire \stat_rd_data[15]_i_2_n_0 ;
  wire \stat_rd_data[15]_i_3_n_0 ;
  wire \stat_rd_data[15]_i_5_n_0 ;
  wire \stat_rd_data[15]_i_6_n_0 ;
  wire \stat_rd_data[15]_i_7_n_0 ;
  wire \stat_rd_data[16]_i_10_n_0 ;
  wire \stat_rd_data[16]_i_11_n_0 ;
  wire \stat_rd_data[16]_i_12_n_0 ;
  wire \stat_rd_data[16]_i_13_n_0 ;
  wire \stat_rd_data[16]_i_14_n_0 ;
  wire \stat_rd_data[16]_i_2_n_0 ;
  wire \stat_rd_data[16]_i_3_n_0 ;
  wire \stat_rd_data[16]_i_5_n_0 ;
  wire \stat_rd_data[16]_i_6_n_0 ;
  wire \stat_rd_data[16]_i_7_n_0 ;
  wire \stat_rd_data[17]_i_10_n_0 ;
  wire \stat_rd_data[17]_i_11_n_0 ;
  wire \stat_rd_data[17]_i_12_n_0 ;
  wire \stat_rd_data[17]_i_13_n_0 ;
  wire \stat_rd_data[17]_i_14_n_0 ;
  wire \stat_rd_data[17]_i_2_n_0 ;
  wire \stat_rd_data[17]_i_3_n_0 ;
  wire \stat_rd_data[17]_i_5_n_0 ;
  wire \stat_rd_data[17]_i_6_n_0 ;
  wire \stat_rd_data[17]_i_7_n_0 ;
  wire \stat_rd_data[18]_i_10_n_0 ;
  wire \stat_rd_data[18]_i_11_n_0 ;
  wire \stat_rd_data[18]_i_12_n_0 ;
  wire \stat_rd_data[18]_i_13_n_0 ;
  wire \stat_rd_data[18]_i_14_n_0 ;
  wire \stat_rd_data[18]_i_2_n_0 ;
  wire \stat_rd_data[18]_i_3_n_0 ;
  wire \stat_rd_data[18]_i_5_n_0 ;
  wire \stat_rd_data[18]_i_6_n_0 ;
  wire \stat_rd_data[18]_i_7_n_0 ;
  wire \stat_rd_data[19]_i_10_n_0 ;
  wire \stat_rd_data[19]_i_11_n_0 ;
  wire \stat_rd_data[19]_i_12_n_0 ;
  wire \stat_rd_data[19]_i_13_n_0 ;
  wire \stat_rd_data[19]_i_14_n_0 ;
  wire \stat_rd_data[19]_i_2_n_0 ;
  wire \stat_rd_data[19]_i_3_n_0 ;
  wire \stat_rd_data[19]_i_5_n_0 ;
  wire \stat_rd_data[19]_i_6_n_0 ;
  wire \stat_rd_data[19]_i_7_n_0 ;
  wire \stat_rd_data[1]_i_10_n_0 ;
  wire \stat_rd_data[1]_i_11_n_0 ;
  wire \stat_rd_data[1]_i_12_n_0 ;
  wire \stat_rd_data[1]_i_13_n_0 ;
  wire \stat_rd_data[1]_i_14_n_0 ;
  wire \stat_rd_data[1]_i_2_n_0 ;
  wire \stat_rd_data[1]_i_3_n_0 ;
  wire \stat_rd_data[1]_i_5_n_0 ;
  wire \stat_rd_data[1]_i_6_n_0 ;
  wire \stat_rd_data[1]_i_7_n_0 ;
  wire \stat_rd_data[20]_i_10_n_0 ;
  wire \stat_rd_data[20]_i_11_n_0 ;
  wire \stat_rd_data[20]_i_12_n_0 ;
  wire \stat_rd_data[20]_i_13_n_0 ;
  wire \stat_rd_data[20]_i_14_n_0 ;
  wire \stat_rd_data[20]_i_2_n_0 ;
  wire \stat_rd_data[20]_i_3_n_0 ;
  wire \stat_rd_data[20]_i_5_n_0 ;
  wire \stat_rd_data[20]_i_6_n_0 ;
  wire \stat_rd_data[20]_i_7_n_0 ;
  wire \stat_rd_data[21]_i_10_n_0 ;
  wire \stat_rd_data[21]_i_11_n_0 ;
  wire \stat_rd_data[21]_i_12_n_0 ;
  wire \stat_rd_data[21]_i_13_n_0 ;
  wire \stat_rd_data[21]_i_14_n_0 ;
  wire \stat_rd_data[21]_i_2_n_0 ;
  wire \stat_rd_data[21]_i_3_n_0 ;
  wire \stat_rd_data[21]_i_5_n_0 ;
  wire \stat_rd_data[21]_i_6_n_0 ;
  wire \stat_rd_data[21]_i_7_n_0 ;
  wire \stat_rd_data[22]_i_10_n_0 ;
  wire \stat_rd_data[22]_i_11_n_0 ;
  wire \stat_rd_data[22]_i_12_n_0 ;
  wire \stat_rd_data[22]_i_13_n_0 ;
  wire \stat_rd_data[22]_i_14_n_0 ;
  wire \stat_rd_data[22]_i_2_n_0 ;
  wire \stat_rd_data[22]_i_3_n_0 ;
  wire \stat_rd_data[22]_i_5_n_0 ;
  wire \stat_rd_data[22]_i_6_n_0 ;
  wire \stat_rd_data[22]_i_7_n_0 ;
  wire \stat_rd_data[23]_i_10_n_0 ;
  wire \stat_rd_data[23]_i_11_n_0 ;
  wire \stat_rd_data[23]_i_12_n_0 ;
  wire \stat_rd_data[23]_i_13_n_0 ;
  wire \stat_rd_data[23]_i_14_n_0 ;
  wire \stat_rd_data[23]_i_2_n_0 ;
  wire \stat_rd_data[23]_i_3_n_0 ;
  wire \stat_rd_data[23]_i_5_n_0 ;
  wire \stat_rd_data[23]_i_6_n_0 ;
  wire \stat_rd_data[23]_i_7_n_0 ;
  wire \stat_rd_data[24]_i_10_n_0 ;
  wire \stat_rd_data[24]_i_11_n_0 ;
  wire \stat_rd_data[24]_i_12_n_0 ;
  wire \stat_rd_data[24]_i_13_n_0 ;
  wire \stat_rd_data[24]_i_14_n_0 ;
  wire \stat_rd_data[24]_i_2_n_0 ;
  wire \stat_rd_data[24]_i_3_n_0 ;
  wire \stat_rd_data[24]_i_5_n_0 ;
  wire \stat_rd_data[24]_i_6_n_0 ;
  wire \stat_rd_data[24]_i_7_n_0 ;
  wire \stat_rd_data[25]_i_10_n_0 ;
  wire \stat_rd_data[25]_i_11_n_0 ;
  wire \stat_rd_data[25]_i_12_n_0 ;
  wire \stat_rd_data[25]_i_13_n_0 ;
  wire \stat_rd_data[25]_i_14_n_0 ;
  wire \stat_rd_data[25]_i_2_n_0 ;
  wire \stat_rd_data[25]_i_3_n_0 ;
  wire \stat_rd_data[25]_i_5_n_0 ;
  wire \stat_rd_data[25]_i_6_n_0 ;
  wire \stat_rd_data[25]_i_7_n_0 ;
  wire \stat_rd_data[26]_i_10_n_0 ;
  wire \stat_rd_data[26]_i_11_n_0 ;
  wire \stat_rd_data[26]_i_12_n_0 ;
  wire \stat_rd_data[26]_i_13_n_0 ;
  wire \stat_rd_data[26]_i_14_n_0 ;
  wire \stat_rd_data[26]_i_2_n_0 ;
  wire \stat_rd_data[26]_i_3_n_0 ;
  wire \stat_rd_data[26]_i_5_n_0 ;
  wire \stat_rd_data[26]_i_6_n_0 ;
  wire \stat_rd_data[26]_i_7_n_0 ;
  wire \stat_rd_data[27]_i_10_n_0 ;
  wire \stat_rd_data[27]_i_11_n_0 ;
  wire \stat_rd_data[27]_i_12_n_0 ;
  wire \stat_rd_data[27]_i_13_n_0 ;
  wire \stat_rd_data[27]_i_14_n_0 ;
  wire \stat_rd_data[27]_i_2_n_0 ;
  wire \stat_rd_data[27]_i_3_n_0 ;
  wire \stat_rd_data[27]_i_5_n_0 ;
  wire \stat_rd_data[27]_i_6_n_0 ;
  wire \stat_rd_data[27]_i_7_n_0 ;
  wire \stat_rd_data[28]_i_10_n_0 ;
  wire \stat_rd_data[28]_i_11_n_0 ;
  wire \stat_rd_data[28]_i_12_n_0 ;
  wire \stat_rd_data[28]_i_13_n_0 ;
  wire \stat_rd_data[28]_i_14_n_0 ;
  wire \stat_rd_data[28]_i_2_n_0 ;
  wire \stat_rd_data[28]_i_3_n_0 ;
  wire \stat_rd_data[28]_i_5_n_0 ;
  wire \stat_rd_data[28]_i_6_n_0 ;
  wire \stat_rd_data[28]_i_7_n_0 ;
  wire \stat_rd_data[29]_i_10_n_0 ;
  wire \stat_rd_data[29]_i_11_n_0 ;
  wire \stat_rd_data[29]_i_12_n_0 ;
  wire \stat_rd_data[29]_i_13_n_0 ;
  wire \stat_rd_data[29]_i_14_n_0 ;
  wire \stat_rd_data[29]_i_2_n_0 ;
  wire \stat_rd_data[29]_i_3_n_0 ;
  wire \stat_rd_data[29]_i_5_n_0 ;
  wire \stat_rd_data[29]_i_6_n_0 ;
  wire \stat_rd_data[29]_i_7_n_0 ;
  wire \stat_rd_data[2]_i_10_n_0 ;
  wire \stat_rd_data[2]_i_11_n_0 ;
  wire \stat_rd_data[2]_i_12_n_0 ;
  wire \stat_rd_data[2]_i_13_n_0 ;
  wire \stat_rd_data[2]_i_14_n_0 ;
  wire \stat_rd_data[2]_i_2_n_0 ;
  wire \stat_rd_data[2]_i_3_n_0 ;
  wire \stat_rd_data[2]_i_5_n_0 ;
  wire \stat_rd_data[2]_i_6_n_0 ;
  wire \stat_rd_data[2]_i_7_n_0 ;
  wire \stat_rd_data[30]_i_10_n_0 ;
  wire \stat_rd_data[30]_i_11_n_0 ;
  wire \stat_rd_data[30]_i_12_n_0 ;
  wire \stat_rd_data[30]_i_13_n_0 ;
  wire \stat_rd_data[30]_i_14_n_0 ;
  wire \stat_rd_data[30]_i_2_n_0 ;
  wire \stat_rd_data[30]_i_3_n_0 ;
  wire \stat_rd_data[30]_i_5_n_0 ;
  wire \stat_rd_data[30]_i_6_n_0 ;
  wire \stat_rd_data[30]_i_7_n_0 ;
  wire \stat_rd_data[31]_i_10_n_0 ;
  wire \stat_rd_data[31]_i_11_n_0 ;
  wire \stat_rd_data[31]_i_12_n_0 ;
  wire \stat_rd_data[31]_i_13_n_0 ;
  wire \stat_rd_data[31]_i_14_n_0 ;
  wire \stat_rd_data[31]_i_2_n_0 ;
  wire \stat_rd_data[31]_i_3_n_0 ;
  wire \stat_rd_data[31]_i_5_n_0 ;
  wire \stat_rd_data[31]_i_6_n_0 ;
  wire \stat_rd_data[31]_i_7_n_0 ;
  wire \stat_rd_data[32]_i_10_n_0 ;
  wire \stat_rd_data[32]_i_11_n_0 ;
  wire \stat_rd_data[32]_i_12_n_0 ;
  wire \stat_rd_data[32]_i_13_n_0 ;
  wire \stat_rd_data[32]_i_14_n_0 ;
  wire \stat_rd_data[32]_i_2_n_0 ;
  wire \stat_rd_data[32]_i_3_n_0 ;
  wire \stat_rd_data[32]_i_5_n_0 ;
  wire \stat_rd_data[32]_i_6_n_0 ;
  wire \stat_rd_data[32]_i_7_n_0 ;
  wire \stat_rd_data[33]_i_10_n_0 ;
  wire \stat_rd_data[33]_i_11_n_0 ;
  wire \stat_rd_data[33]_i_12_n_0 ;
  wire \stat_rd_data[33]_i_13_n_0 ;
  wire \stat_rd_data[33]_i_14_n_0 ;
  wire \stat_rd_data[33]_i_2_n_0 ;
  wire \stat_rd_data[33]_i_3_n_0 ;
  wire \stat_rd_data[33]_i_5_n_0 ;
  wire \stat_rd_data[33]_i_6_n_0 ;
  wire \stat_rd_data[33]_i_7_n_0 ;
  wire \stat_rd_data[34]_i_10_n_0 ;
  wire \stat_rd_data[34]_i_11_n_0 ;
  wire \stat_rd_data[34]_i_12_n_0 ;
  wire \stat_rd_data[34]_i_13_n_0 ;
  wire \stat_rd_data[34]_i_14_n_0 ;
  wire \stat_rd_data[34]_i_2_n_0 ;
  wire \stat_rd_data[34]_i_3_n_0 ;
  wire \stat_rd_data[34]_i_5_n_0 ;
  wire \stat_rd_data[34]_i_6_n_0 ;
  wire \stat_rd_data[34]_i_7_n_0 ;
  wire \stat_rd_data[35]_i_10_n_0 ;
  wire \stat_rd_data[35]_i_11_n_0 ;
  wire \stat_rd_data[35]_i_12_n_0 ;
  wire \stat_rd_data[35]_i_13_n_0 ;
  wire \stat_rd_data[35]_i_14_n_0 ;
  wire \stat_rd_data[35]_i_2_n_0 ;
  wire \stat_rd_data[35]_i_3_n_0 ;
  wire \stat_rd_data[35]_i_5_n_0 ;
  wire \stat_rd_data[35]_i_6_n_0 ;
  wire \stat_rd_data[35]_i_7_n_0 ;
  wire \stat_rd_data[36]_i_10_n_0 ;
  wire \stat_rd_data[36]_i_11_n_0 ;
  wire \stat_rd_data[36]_i_12_n_0 ;
  wire \stat_rd_data[36]_i_13_n_0 ;
  wire \stat_rd_data[36]_i_14_n_0 ;
  wire \stat_rd_data[36]_i_2_n_0 ;
  wire \stat_rd_data[36]_i_3_n_0 ;
  wire \stat_rd_data[36]_i_5_n_0 ;
  wire \stat_rd_data[36]_i_6_n_0 ;
  wire \stat_rd_data[36]_i_7_n_0 ;
  wire \stat_rd_data[37]_i_10_n_0 ;
  wire \stat_rd_data[37]_i_11_n_0 ;
  wire \stat_rd_data[37]_i_12_n_0 ;
  wire \stat_rd_data[37]_i_13_n_0 ;
  wire \stat_rd_data[37]_i_14_n_0 ;
  wire \stat_rd_data[37]_i_2_n_0 ;
  wire \stat_rd_data[37]_i_3_n_0 ;
  wire \stat_rd_data[37]_i_5_n_0 ;
  wire \stat_rd_data[37]_i_6_n_0 ;
  wire \stat_rd_data[37]_i_7_n_0 ;
  wire \stat_rd_data[38]_i_10_n_0 ;
  wire \stat_rd_data[38]_i_11_n_0 ;
  wire \stat_rd_data[38]_i_12_n_0 ;
  wire \stat_rd_data[38]_i_13_n_0 ;
  wire \stat_rd_data[38]_i_14_n_0 ;
  wire \stat_rd_data[38]_i_2_n_0 ;
  wire \stat_rd_data[38]_i_3_n_0 ;
  wire \stat_rd_data[38]_i_5_n_0 ;
  wire \stat_rd_data[38]_i_6_n_0 ;
  wire \stat_rd_data[38]_i_7_n_0 ;
  wire \stat_rd_data[39]_i_10_n_0 ;
  wire \stat_rd_data[39]_i_11_n_0 ;
  wire \stat_rd_data[39]_i_12_n_0 ;
  wire \stat_rd_data[39]_i_13_n_0 ;
  wire \stat_rd_data[39]_i_14_n_0 ;
  wire \stat_rd_data[39]_i_2_n_0 ;
  wire \stat_rd_data[39]_i_3_n_0 ;
  wire \stat_rd_data[39]_i_5_n_0 ;
  wire \stat_rd_data[39]_i_6_n_0 ;
  wire \stat_rd_data[39]_i_7_n_0 ;
  wire \stat_rd_data[3]_i_10_n_0 ;
  wire \stat_rd_data[3]_i_11_n_0 ;
  wire \stat_rd_data[3]_i_12_n_0 ;
  wire \stat_rd_data[3]_i_13_n_0 ;
  wire \stat_rd_data[3]_i_14_n_0 ;
  wire \stat_rd_data[3]_i_2_n_0 ;
  wire \stat_rd_data[3]_i_3_n_0 ;
  wire \stat_rd_data[3]_i_5_n_0 ;
  wire \stat_rd_data[3]_i_6_n_0 ;
  wire \stat_rd_data[3]_i_7_n_0 ;
  wire \stat_rd_data[40]_i_10_n_0 ;
  wire \stat_rd_data[40]_i_11_n_0 ;
  wire \stat_rd_data[40]_i_12_n_0 ;
  wire \stat_rd_data[40]_i_13_n_0 ;
  wire \stat_rd_data[40]_i_14_n_0 ;
  wire \stat_rd_data[40]_i_2_n_0 ;
  wire \stat_rd_data[40]_i_3_n_0 ;
  wire \stat_rd_data[40]_i_5_n_0 ;
  wire \stat_rd_data[40]_i_6_n_0 ;
  wire \stat_rd_data[40]_i_7_n_0 ;
  wire \stat_rd_data[41]_i_10_n_0 ;
  wire \stat_rd_data[41]_i_11_n_0 ;
  wire \stat_rd_data[41]_i_12_n_0 ;
  wire \stat_rd_data[41]_i_13_n_0 ;
  wire \stat_rd_data[41]_i_14_n_0 ;
  wire \stat_rd_data[41]_i_2_n_0 ;
  wire \stat_rd_data[41]_i_3_n_0 ;
  wire \stat_rd_data[41]_i_5_n_0 ;
  wire \stat_rd_data[41]_i_6_n_0 ;
  wire \stat_rd_data[41]_i_7_n_0 ;
  wire \stat_rd_data[42]_i_10_n_0 ;
  wire \stat_rd_data[42]_i_11_n_0 ;
  wire \stat_rd_data[42]_i_12_n_0 ;
  wire \stat_rd_data[42]_i_13_n_0 ;
  wire \stat_rd_data[42]_i_14_n_0 ;
  wire \stat_rd_data[42]_i_2_n_0 ;
  wire \stat_rd_data[42]_i_3_n_0 ;
  wire \stat_rd_data[42]_i_5_n_0 ;
  wire \stat_rd_data[42]_i_6_n_0 ;
  wire \stat_rd_data[42]_i_7_n_0 ;
  wire \stat_rd_data[43]_i_10_n_0 ;
  wire \stat_rd_data[43]_i_11_n_0 ;
  wire \stat_rd_data[43]_i_12_n_0 ;
  wire \stat_rd_data[43]_i_13_n_0 ;
  wire \stat_rd_data[43]_i_14_n_0 ;
  wire \stat_rd_data[43]_i_2_n_0 ;
  wire \stat_rd_data[43]_i_3_n_0 ;
  wire \stat_rd_data[43]_i_5_n_0 ;
  wire \stat_rd_data[43]_i_6_n_0 ;
  wire \stat_rd_data[43]_i_7_n_0 ;
  wire \stat_rd_data[44]_i_10_n_0 ;
  wire \stat_rd_data[44]_i_11_n_0 ;
  wire \stat_rd_data[44]_i_12_n_0 ;
  wire \stat_rd_data[44]_i_13_n_0 ;
  wire \stat_rd_data[44]_i_14_n_0 ;
  wire \stat_rd_data[44]_i_2_n_0 ;
  wire \stat_rd_data[44]_i_3_n_0 ;
  wire \stat_rd_data[44]_i_5_n_0 ;
  wire \stat_rd_data[44]_i_6_n_0 ;
  wire \stat_rd_data[44]_i_7_n_0 ;
  wire \stat_rd_data[45]_i_10_n_0 ;
  wire \stat_rd_data[45]_i_11_n_0 ;
  wire \stat_rd_data[45]_i_12_n_0 ;
  wire \stat_rd_data[45]_i_13_n_0 ;
  wire \stat_rd_data[45]_i_14_n_0 ;
  wire \stat_rd_data[45]_i_2_n_0 ;
  wire \stat_rd_data[45]_i_3_n_0 ;
  wire \stat_rd_data[45]_i_5_n_0 ;
  wire \stat_rd_data[45]_i_6_n_0 ;
  wire \stat_rd_data[45]_i_7_n_0 ;
  wire \stat_rd_data[46]_i_10_n_0 ;
  wire \stat_rd_data[46]_i_11_n_0 ;
  wire \stat_rd_data[46]_i_12_n_0 ;
  wire \stat_rd_data[46]_i_13_n_0 ;
  wire \stat_rd_data[46]_i_14_n_0 ;
  wire \stat_rd_data[46]_i_2_n_0 ;
  wire \stat_rd_data[46]_i_3_n_0 ;
  wire \stat_rd_data[46]_i_5_n_0 ;
  wire \stat_rd_data[46]_i_6_n_0 ;
  wire \stat_rd_data[46]_i_7_n_0 ;
  wire \stat_rd_data[47]_i_10_n_0 ;
  wire \stat_rd_data[47]_i_11_n_0 ;
  wire \stat_rd_data[47]_i_12_n_0 ;
  wire \stat_rd_data[47]_i_13_n_0 ;
  wire \stat_rd_data[47]_i_14_n_0 ;
  wire \stat_rd_data[47]_i_2_n_0 ;
  wire \stat_rd_data[47]_i_3_n_0 ;
  wire \stat_rd_data[47]_i_5_n_0 ;
  wire \stat_rd_data[47]_i_6_n_0 ;
  wire \stat_rd_data[47]_i_7_n_0 ;
  wire \stat_rd_data[48]_i_10_n_0 ;
  wire \stat_rd_data[48]_i_11_n_0 ;
  wire \stat_rd_data[48]_i_12_n_0 ;
  wire \stat_rd_data[48]_i_13_n_0 ;
  wire \stat_rd_data[48]_i_14_n_0 ;
  wire \stat_rd_data[48]_i_2_n_0 ;
  wire \stat_rd_data[48]_i_3_n_0 ;
  wire \stat_rd_data[48]_i_5_n_0 ;
  wire \stat_rd_data[48]_i_6_n_0 ;
  wire \stat_rd_data[48]_i_7_n_0 ;
  wire \stat_rd_data[49]_i_10_n_0 ;
  wire \stat_rd_data[49]_i_11_n_0 ;
  wire \stat_rd_data[49]_i_12_n_0 ;
  wire \stat_rd_data[49]_i_13_n_0 ;
  wire \stat_rd_data[49]_i_14_n_0 ;
  wire \stat_rd_data[49]_i_2_n_0 ;
  wire \stat_rd_data[49]_i_3_n_0 ;
  wire \stat_rd_data[49]_i_5_n_0 ;
  wire \stat_rd_data[49]_i_6_n_0 ;
  wire \stat_rd_data[49]_i_7_n_0 ;
  wire \stat_rd_data[4]_i_10_n_0 ;
  wire \stat_rd_data[4]_i_11_n_0 ;
  wire \stat_rd_data[4]_i_12_n_0 ;
  wire \stat_rd_data[4]_i_13_n_0 ;
  wire \stat_rd_data[4]_i_14_n_0 ;
  wire \stat_rd_data[4]_i_2_n_0 ;
  wire \stat_rd_data[4]_i_3_n_0 ;
  wire \stat_rd_data[4]_i_5_n_0 ;
  wire \stat_rd_data[4]_i_6_n_0 ;
  wire \stat_rd_data[4]_i_7_n_0 ;
  wire \stat_rd_data[50]_i_10_n_0 ;
  wire \stat_rd_data[50]_i_11_n_0 ;
  wire \stat_rd_data[50]_i_12_n_0 ;
  wire \stat_rd_data[50]_i_13_n_0 ;
  wire \stat_rd_data[50]_i_14_n_0 ;
  wire \stat_rd_data[50]_i_2_n_0 ;
  wire \stat_rd_data[50]_i_3_n_0 ;
  wire \stat_rd_data[50]_i_5_n_0 ;
  wire \stat_rd_data[50]_i_6_n_0 ;
  wire \stat_rd_data[50]_i_7_n_0 ;
  wire \stat_rd_data[51]_i_10_n_0 ;
  wire \stat_rd_data[51]_i_11_n_0 ;
  wire \stat_rd_data[51]_i_12_n_0 ;
  wire \stat_rd_data[51]_i_13_n_0 ;
  wire \stat_rd_data[51]_i_14_n_0 ;
  wire \stat_rd_data[51]_i_2_n_0 ;
  wire \stat_rd_data[51]_i_3_n_0 ;
  wire \stat_rd_data[51]_i_5_n_0 ;
  wire \stat_rd_data[51]_i_6_n_0 ;
  wire \stat_rd_data[51]_i_7_n_0 ;
  wire \stat_rd_data[52]_i_10_n_0 ;
  wire \stat_rd_data[52]_i_11_n_0 ;
  wire \stat_rd_data[52]_i_12_n_0 ;
  wire \stat_rd_data[52]_i_13_n_0 ;
  wire \stat_rd_data[52]_i_14_n_0 ;
  wire \stat_rd_data[52]_i_2_n_0 ;
  wire \stat_rd_data[52]_i_3_n_0 ;
  wire \stat_rd_data[52]_i_5_n_0 ;
  wire \stat_rd_data[52]_i_6_n_0 ;
  wire \stat_rd_data[52]_i_7_n_0 ;
  wire \stat_rd_data[53]_i_10_n_0 ;
  wire \stat_rd_data[53]_i_11_n_0 ;
  wire \stat_rd_data[53]_i_12_n_0 ;
  wire \stat_rd_data[53]_i_13_n_0 ;
  wire \stat_rd_data[53]_i_14_n_0 ;
  wire \stat_rd_data[53]_i_2_n_0 ;
  wire \stat_rd_data[53]_i_3_n_0 ;
  wire \stat_rd_data[53]_i_5_n_0 ;
  wire \stat_rd_data[53]_i_6_n_0 ;
  wire \stat_rd_data[53]_i_7_n_0 ;
  wire \stat_rd_data[54]_i_10_n_0 ;
  wire \stat_rd_data[54]_i_11_n_0 ;
  wire \stat_rd_data[54]_i_12_n_0 ;
  wire \stat_rd_data[54]_i_13_n_0 ;
  wire \stat_rd_data[54]_i_14_n_0 ;
  wire \stat_rd_data[54]_i_2_n_0 ;
  wire \stat_rd_data[54]_i_3_n_0 ;
  wire \stat_rd_data[54]_i_5_n_0 ;
  wire \stat_rd_data[54]_i_6_n_0 ;
  wire \stat_rd_data[54]_i_7_n_0 ;
  wire \stat_rd_data[55]_i_10_n_0 ;
  wire \stat_rd_data[55]_i_11_n_0 ;
  wire \stat_rd_data[55]_i_12_n_0 ;
  wire \stat_rd_data[55]_i_13_n_0 ;
  wire \stat_rd_data[55]_i_14_n_0 ;
  wire \stat_rd_data[55]_i_2_n_0 ;
  wire \stat_rd_data[55]_i_3_n_0 ;
  wire \stat_rd_data[55]_i_5_n_0 ;
  wire \stat_rd_data[55]_i_6_n_0 ;
  wire \stat_rd_data[55]_i_7_n_0 ;
  wire \stat_rd_data[56]_i_10_n_0 ;
  wire \stat_rd_data[56]_i_11_n_0 ;
  wire \stat_rd_data[56]_i_12_n_0 ;
  wire \stat_rd_data[56]_i_13_n_0 ;
  wire \stat_rd_data[56]_i_14_n_0 ;
  wire \stat_rd_data[56]_i_2_n_0 ;
  wire \stat_rd_data[56]_i_3_n_0 ;
  wire \stat_rd_data[56]_i_5_n_0 ;
  wire \stat_rd_data[56]_i_6_n_0 ;
  wire \stat_rd_data[56]_i_7_n_0 ;
  wire \stat_rd_data[57]_i_10_n_0 ;
  wire \stat_rd_data[57]_i_11_n_0 ;
  wire \stat_rd_data[57]_i_12_n_0 ;
  wire \stat_rd_data[57]_i_13_n_0 ;
  wire \stat_rd_data[57]_i_14_n_0 ;
  wire \stat_rd_data[57]_i_2_n_0 ;
  wire \stat_rd_data[57]_i_3_n_0 ;
  wire \stat_rd_data[57]_i_5_n_0 ;
  wire \stat_rd_data[57]_i_6_n_0 ;
  wire \stat_rd_data[57]_i_7_n_0 ;
  wire \stat_rd_data[58]_i_10_n_0 ;
  wire \stat_rd_data[58]_i_11_n_0 ;
  wire \stat_rd_data[58]_i_12_n_0 ;
  wire \stat_rd_data[58]_i_13_n_0 ;
  wire \stat_rd_data[58]_i_14_n_0 ;
  wire \stat_rd_data[58]_i_2_n_0 ;
  wire \stat_rd_data[58]_i_3_n_0 ;
  wire \stat_rd_data[58]_i_5_n_0 ;
  wire \stat_rd_data[58]_i_6_n_0 ;
  wire \stat_rd_data[58]_i_7_n_0 ;
  wire \stat_rd_data[59]_i_10_n_0 ;
  wire \stat_rd_data[59]_i_11_n_0 ;
  wire \stat_rd_data[59]_i_12_n_0 ;
  wire \stat_rd_data[59]_i_13_n_0 ;
  wire \stat_rd_data[59]_i_14_n_0 ;
  wire \stat_rd_data[59]_i_2_n_0 ;
  wire \stat_rd_data[59]_i_3_n_0 ;
  wire \stat_rd_data[59]_i_5_n_0 ;
  wire \stat_rd_data[59]_i_6_n_0 ;
  wire \stat_rd_data[59]_i_7_n_0 ;
  wire \stat_rd_data[5]_i_10_n_0 ;
  wire \stat_rd_data[5]_i_11_n_0 ;
  wire \stat_rd_data[5]_i_12_n_0 ;
  wire \stat_rd_data[5]_i_13_n_0 ;
  wire \stat_rd_data[5]_i_14_n_0 ;
  wire \stat_rd_data[5]_i_2_n_0 ;
  wire \stat_rd_data[5]_i_3_n_0 ;
  wire \stat_rd_data[5]_i_5_n_0 ;
  wire \stat_rd_data[5]_i_6_n_0 ;
  wire \stat_rd_data[5]_i_7_n_0 ;
  wire \stat_rd_data[60]_i_10_n_0 ;
  wire \stat_rd_data[60]_i_11_n_0 ;
  wire \stat_rd_data[60]_i_12_n_0 ;
  wire \stat_rd_data[60]_i_13_n_0 ;
  wire \stat_rd_data[60]_i_14_n_0 ;
  wire \stat_rd_data[60]_i_2_n_0 ;
  wire \stat_rd_data[60]_i_3_n_0 ;
  wire \stat_rd_data[60]_i_5_n_0 ;
  wire \stat_rd_data[60]_i_6_n_0 ;
  wire \stat_rd_data[60]_i_7_n_0 ;
  wire \stat_rd_data[61]_i_10_n_0 ;
  wire \stat_rd_data[61]_i_11_n_0 ;
  wire \stat_rd_data[61]_i_12_n_0 ;
  wire \stat_rd_data[61]_i_13_n_0 ;
  wire \stat_rd_data[61]_i_14_n_0 ;
  wire \stat_rd_data[61]_i_2_n_0 ;
  wire \stat_rd_data[61]_i_3_n_0 ;
  wire \stat_rd_data[61]_i_5_n_0 ;
  wire \stat_rd_data[61]_i_6_n_0 ;
  wire \stat_rd_data[61]_i_7_n_0 ;
  wire \stat_rd_data[62]_i_10_n_0 ;
  wire \stat_rd_data[62]_i_11_n_0 ;
  wire \stat_rd_data[62]_i_12_n_0 ;
  wire \stat_rd_data[62]_i_13_n_0 ;
  wire \stat_rd_data[62]_i_14_n_0 ;
  wire \stat_rd_data[62]_i_2_n_0 ;
  wire \stat_rd_data[62]_i_3_n_0 ;
  wire \stat_rd_data[62]_i_5_n_0 ;
  wire \stat_rd_data[62]_i_6_n_0 ;
  wire \stat_rd_data[62]_i_7_n_0 ;
  wire \stat_rd_data[63]_i_10_n_0 ;
  wire \stat_rd_data[63]_i_11_n_0 ;
  wire \stat_rd_data[63]_i_12_n_0 ;
  wire \stat_rd_data[63]_i_13_n_0 ;
  wire \stat_rd_data[63]_i_16_n_0 ;
  wire \stat_rd_data[63]_i_17_n_0 ;
  wire \stat_rd_data[63]_i_18_n_0 ;
  wire \stat_rd_data[63]_i_19_n_0 ;
  wire \stat_rd_data[63]_i_1_n_0 ;
  wire \stat_rd_data[63]_i_20_n_0 ;
  wire \stat_rd_data[63]_i_3_n_0 ;
  wire \stat_rd_data[63]_i_4_n_0 ;
  wire \stat_rd_data[63]_i_5_n_0 ;
  wire \stat_rd_data[63]_i_6_n_0 ;
  wire \stat_rd_data[63]_i_7_n_0 ;
  wire \stat_rd_data[63]_i_9_n_0 ;
  wire \stat_rd_data[6]_i_10_n_0 ;
  wire \stat_rd_data[6]_i_11_n_0 ;
  wire \stat_rd_data[6]_i_12_n_0 ;
  wire \stat_rd_data[6]_i_13_n_0 ;
  wire \stat_rd_data[6]_i_14_n_0 ;
  wire \stat_rd_data[6]_i_2_n_0 ;
  wire \stat_rd_data[6]_i_3_n_0 ;
  wire \stat_rd_data[6]_i_5_n_0 ;
  wire \stat_rd_data[6]_i_6_n_0 ;
  wire \stat_rd_data[6]_i_7_n_0 ;
  wire \stat_rd_data[7]_i_10_n_0 ;
  wire \stat_rd_data[7]_i_11_n_0 ;
  wire \stat_rd_data[7]_i_12_n_0 ;
  wire \stat_rd_data[7]_i_13_n_0 ;
  wire \stat_rd_data[7]_i_14_n_0 ;
  wire \stat_rd_data[7]_i_2_n_0 ;
  wire \stat_rd_data[7]_i_3_n_0 ;
  wire \stat_rd_data[7]_i_5_n_0 ;
  wire \stat_rd_data[7]_i_6_n_0 ;
  wire \stat_rd_data[7]_i_7_n_0 ;
  wire \stat_rd_data[8]_i_10_n_0 ;
  wire \stat_rd_data[8]_i_11_n_0 ;
  wire \stat_rd_data[8]_i_12_n_0 ;
  wire \stat_rd_data[8]_i_13_n_0 ;
  wire \stat_rd_data[8]_i_14_n_0 ;
  wire \stat_rd_data[8]_i_2_n_0 ;
  wire \stat_rd_data[8]_i_3_n_0 ;
  wire \stat_rd_data[8]_i_5_n_0 ;
  wire \stat_rd_data[8]_i_6_n_0 ;
  wire \stat_rd_data[8]_i_7_n_0 ;
  wire \stat_rd_data[9]_i_10_n_0 ;
  wire \stat_rd_data[9]_i_11_n_0 ;
  wire \stat_rd_data[9]_i_12_n_0 ;
  wire \stat_rd_data[9]_i_13_n_0 ;
  wire \stat_rd_data[9]_i_14_n_0 ;
  wire \stat_rd_data[9]_i_2_n_0 ;
  wire \stat_rd_data[9]_i_3_n_0 ;
  wire \stat_rd_data[9]_i_5_n_0 ;
  wire \stat_rd_data[9]_i_6_n_0 ;
  wire \stat_rd_data[9]_i_7_n_0 ;
  wire \stat_rd_data_reg[0]_i_4_n_0 ;
  wire \stat_rd_data_reg[0]_i_8_n_0 ;
  wire \stat_rd_data_reg[0]_i_9_n_0 ;
  wire \stat_rd_data_reg[10]_i_4_n_0 ;
  wire \stat_rd_data_reg[10]_i_8_n_0 ;
  wire \stat_rd_data_reg[10]_i_9_n_0 ;
  wire \stat_rd_data_reg[11]_i_4_n_0 ;
  wire \stat_rd_data_reg[11]_i_8_n_0 ;
  wire \stat_rd_data_reg[11]_i_9_n_0 ;
  wire \stat_rd_data_reg[12]_i_4_n_0 ;
  wire \stat_rd_data_reg[12]_i_8_n_0 ;
  wire \stat_rd_data_reg[12]_i_9_n_0 ;
  wire \stat_rd_data_reg[13]_i_4_n_0 ;
  wire \stat_rd_data_reg[13]_i_8_n_0 ;
  wire \stat_rd_data_reg[13]_i_9_n_0 ;
  wire \stat_rd_data_reg[14]_i_4_n_0 ;
  wire \stat_rd_data_reg[14]_i_8_n_0 ;
  wire \stat_rd_data_reg[14]_i_9_n_0 ;
  wire \stat_rd_data_reg[15]_i_4_n_0 ;
  wire \stat_rd_data_reg[15]_i_8_n_0 ;
  wire \stat_rd_data_reg[15]_i_9_n_0 ;
  wire \stat_rd_data_reg[16]_i_4_n_0 ;
  wire \stat_rd_data_reg[16]_i_8_n_0 ;
  wire \stat_rd_data_reg[16]_i_9_n_0 ;
  wire \stat_rd_data_reg[17]_i_4_n_0 ;
  wire \stat_rd_data_reg[17]_i_8_n_0 ;
  wire \stat_rd_data_reg[17]_i_9_n_0 ;
  wire \stat_rd_data_reg[18]_i_4_n_0 ;
  wire \stat_rd_data_reg[18]_i_8_n_0 ;
  wire \stat_rd_data_reg[18]_i_9_n_0 ;
  wire \stat_rd_data_reg[19]_i_4_n_0 ;
  wire \stat_rd_data_reg[19]_i_8_n_0 ;
  wire \stat_rd_data_reg[19]_i_9_n_0 ;
  wire \stat_rd_data_reg[1]_i_4_n_0 ;
  wire \stat_rd_data_reg[1]_i_8_n_0 ;
  wire \stat_rd_data_reg[1]_i_9_n_0 ;
  wire \stat_rd_data_reg[20]_i_4_n_0 ;
  wire \stat_rd_data_reg[20]_i_8_n_0 ;
  wire \stat_rd_data_reg[20]_i_9_n_0 ;
  wire \stat_rd_data_reg[21]_i_4_n_0 ;
  wire \stat_rd_data_reg[21]_i_8_n_0 ;
  wire \stat_rd_data_reg[21]_i_9_n_0 ;
  wire \stat_rd_data_reg[22]_i_4_n_0 ;
  wire \stat_rd_data_reg[22]_i_8_n_0 ;
  wire \stat_rd_data_reg[22]_i_9_n_0 ;
  wire \stat_rd_data_reg[23]_i_4_n_0 ;
  wire \stat_rd_data_reg[23]_i_8_n_0 ;
  wire \stat_rd_data_reg[23]_i_9_n_0 ;
  wire \stat_rd_data_reg[24]_i_4_n_0 ;
  wire \stat_rd_data_reg[24]_i_8_n_0 ;
  wire \stat_rd_data_reg[24]_i_9_n_0 ;
  wire \stat_rd_data_reg[25]_i_4_n_0 ;
  wire \stat_rd_data_reg[25]_i_8_n_0 ;
  wire \stat_rd_data_reg[25]_i_9_n_0 ;
  wire \stat_rd_data_reg[26]_i_4_n_0 ;
  wire \stat_rd_data_reg[26]_i_8_n_0 ;
  wire \stat_rd_data_reg[26]_i_9_n_0 ;
  wire \stat_rd_data_reg[27]_i_4_n_0 ;
  wire \stat_rd_data_reg[27]_i_8_n_0 ;
  wire \stat_rd_data_reg[27]_i_9_n_0 ;
  wire \stat_rd_data_reg[28]_i_4_n_0 ;
  wire \stat_rd_data_reg[28]_i_8_n_0 ;
  wire \stat_rd_data_reg[28]_i_9_n_0 ;
  wire \stat_rd_data_reg[29]_i_4_n_0 ;
  wire \stat_rd_data_reg[29]_i_8_n_0 ;
  wire \stat_rd_data_reg[29]_i_9_n_0 ;
  wire \stat_rd_data_reg[2]_i_4_n_0 ;
  wire \stat_rd_data_reg[2]_i_8_n_0 ;
  wire \stat_rd_data_reg[2]_i_9_n_0 ;
  wire \stat_rd_data_reg[30]_i_4_n_0 ;
  wire \stat_rd_data_reg[30]_i_8_n_0 ;
  wire \stat_rd_data_reg[30]_i_9_n_0 ;
  wire \stat_rd_data_reg[31]_i_4_n_0 ;
  wire \stat_rd_data_reg[31]_i_8_n_0 ;
  wire \stat_rd_data_reg[31]_i_9_n_0 ;
  wire \stat_rd_data_reg[32]_i_4_n_0 ;
  wire \stat_rd_data_reg[32]_i_8_n_0 ;
  wire \stat_rd_data_reg[32]_i_9_n_0 ;
  wire \stat_rd_data_reg[33]_i_4_n_0 ;
  wire \stat_rd_data_reg[33]_i_8_n_0 ;
  wire \stat_rd_data_reg[33]_i_9_n_0 ;
  wire \stat_rd_data_reg[34]_i_4_n_0 ;
  wire \stat_rd_data_reg[34]_i_8_n_0 ;
  wire \stat_rd_data_reg[34]_i_9_n_0 ;
  wire \stat_rd_data_reg[35]_i_4_n_0 ;
  wire \stat_rd_data_reg[35]_i_8_n_0 ;
  wire \stat_rd_data_reg[35]_i_9_n_0 ;
  wire \stat_rd_data_reg[36]_i_4_n_0 ;
  wire \stat_rd_data_reg[36]_i_8_n_0 ;
  wire \stat_rd_data_reg[36]_i_9_n_0 ;
  wire \stat_rd_data_reg[37]_i_4_n_0 ;
  wire \stat_rd_data_reg[37]_i_8_n_0 ;
  wire \stat_rd_data_reg[37]_i_9_n_0 ;
  wire \stat_rd_data_reg[38]_i_4_n_0 ;
  wire \stat_rd_data_reg[38]_i_8_n_0 ;
  wire \stat_rd_data_reg[38]_i_9_n_0 ;
  wire \stat_rd_data_reg[39]_i_4_n_0 ;
  wire \stat_rd_data_reg[39]_i_8_n_0 ;
  wire \stat_rd_data_reg[39]_i_9_n_0 ;
  wire \stat_rd_data_reg[3]_i_4_n_0 ;
  wire \stat_rd_data_reg[3]_i_8_n_0 ;
  wire \stat_rd_data_reg[3]_i_9_n_0 ;
  wire \stat_rd_data_reg[40]_i_4_n_0 ;
  wire \stat_rd_data_reg[40]_i_8_n_0 ;
  wire \stat_rd_data_reg[40]_i_9_n_0 ;
  wire \stat_rd_data_reg[41]_i_4_n_0 ;
  wire \stat_rd_data_reg[41]_i_8_n_0 ;
  wire \stat_rd_data_reg[41]_i_9_n_0 ;
  wire \stat_rd_data_reg[42]_i_4_n_0 ;
  wire \stat_rd_data_reg[42]_i_8_n_0 ;
  wire \stat_rd_data_reg[42]_i_9_n_0 ;
  wire \stat_rd_data_reg[43]_i_4_n_0 ;
  wire \stat_rd_data_reg[43]_i_8_n_0 ;
  wire \stat_rd_data_reg[43]_i_9_n_0 ;
  wire \stat_rd_data_reg[44]_i_4_n_0 ;
  wire \stat_rd_data_reg[44]_i_8_n_0 ;
  wire \stat_rd_data_reg[44]_i_9_n_0 ;
  wire \stat_rd_data_reg[45]_i_4_n_0 ;
  wire \stat_rd_data_reg[45]_i_8_n_0 ;
  wire \stat_rd_data_reg[45]_i_9_n_0 ;
  wire \stat_rd_data_reg[46]_i_4_n_0 ;
  wire \stat_rd_data_reg[46]_i_8_n_0 ;
  wire \stat_rd_data_reg[46]_i_9_n_0 ;
  wire \stat_rd_data_reg[47]_i_4_n_0 ;
  wire \stat_rd_data_reg[47]_i_8_n_0 ;
  wire \stat_rd_data_reg[47]_i_9_n_0 ;
  wire \stat_rd_data_reg[48]_i_4_n_0 ;
  wire \stat_rd_data_reg[48]_i_8_n_0 ;
  wire \stat_rd_data_reg[48]_i_9_n_0 ;
  wire \stat_rd_data_reg[49]_i_4_n_0 ;
  wire \stat_rd_data_reg[49]_i_8_n_0 ;
  wire \stat_rd_data_reg[49]_i_9_n_0 ;
  wire \stat_rd_data_reg[4]_i_4_n_0 ;
  wire \stat_rd_data_reg[4]_i_8_n_0 ;
  wire \stat_rd_data_reg[4]_i_9_n_0 ;
  wire \stat_rd_data_reg[50]_i_4_n_0 ;
  wire \stat_rd_data_reg[50]_i_8_n_0 ;
  wire \stat_rd_data_reg[50]_i_9_n_0 ;
  wire \stat_rd_data_reg[51]_i_4_n_0 ;
  wire \stat_rd_data_reg[51]_i_8_n_0 ;
  wire \stat_rd_data_reg[51]_i_9_n_0 ;
  wire \stat_rd_data_reg[52]_i_4_n_0 ;
  wire \stat_rd_data_reg[52]_i_8_n_0 ;
  wire \stat_rd_data_reg[52]_i_9_n_0 ;
  wire \stat_rd_data_reg[53]_i_4_n_0 ;
  wire \stat_rd_data_reg[53]_i_8_n_0 ;
  wire \stat_rd_data_reg[53]_i_9_n_0 ;
  wire \stat_rd_data_reg[54]_i_4_n_0 ;
  wire \stat_rd_data_reg[54]_i_8_n_0 ;
  wire \stat_rd_data_reg[54]_i_9_n_0 ;
  wire \stat_rd_data_reg[55]_i_4_n_0 ;
  wire \stat_rd_data_reg[55]_i_8_n_0 ;
  wire \stat_rd_data_reg[55]_i_9_n_0 ;
  wire \stat_rd_data_reg[56]_i_4_n_0 ;
  wire \stat_rd_data_reg[56]_i_8_n_0 ;
  wire \stat_rd_data_reg[56]_i_9_n_0 ;
  wire \stat_rd_data_reg[57]_i_4_n_0 ;
  wire \stat_rd_data_reg[57]_i_8_n_0 ;
  wire \stat_rd_data_reg[57]_i_9_n_0 ;
  wire \stat_rd_data_reg[58]_i_4_n_0 ;
  wire \stat_rd_data_reg[58]_i_8_n_0 ;
  wire \stat_rd_data_reg[58]_i_9_n_0 ;
  wire \stat_rd_data_reg[59]_i_4_n_0 ;
  wire \stat_rd_data_reg[59]_i_8_n_0 ;
  wire \stat_rd_data_reg[59]_i_9_n_0 ;
  wire \stat_rd_data_reg[5]_i_4_n_0 ;
  wire \stat_rd_data_reg[5]_i_8_n_0 ;
  wire \stat_rd_data_reg[5]_i_9_n_0 ;
  wire \stat_rd_data_reg[60]_i_4_n_0 ;
  wire \stat_rd_data_reg[60]_i_8_n_0 ;
  wire \stat_rd_data_reg[60]_i_9_n_0 ;
  wire \stat_rd_data_reg[61]_i_4_n_0 ;
  wire \stat_rd_data_reg[61]_i_8_n_0 ;
  wire \stat_rd_data_reg[61]_i_9_n_0 ;
  wire \stat_rd_data_reg[62]_i_4_n_0 ;
  wire \stat_rd_data_reg[62]_i_8_n_0 ;
  wire \stat_rd_data_reg[62]_i_9_n_0 ;
  wire \stat_rd_data_reg[63]_0 ;
  wire \stat_rd_data_reg[63]_1 ;
  wire \stat_rd_data_reg[63]_i_14_n_0 ;
  wire \stat_rd_data_reg[63]_i_15_n_0 ;
  wire \stat_rd_data_reg[63]_i_8_n_0 ;
  wire \stat_rd_data_reg[6]_i_4_n_0 ;
  wire \stat_rd_data_reg[6]_i_8_n_0 ;
  wire \stat_rd_data_reg[6]_i_9_n_0 ;
  wire \stat_rd_data_reg[7]_i_4_n_0 ;
  wire \stat_rd_data_reg[7]_i_8_n_0 ;
  wire \stat_rd_data_reg[7]_i_9_n_0 ;
  wire \stat_rd_data_reg[8]_i_4_n_0 ;
  wire \stat_rd_data_reg[8]_i_8_n_0 ;
  wire \stat_rd_data_reg[8]_i_9_n_0 ;
  wire \stat_rd_data_reg[9]_i_4_n_0 ;
  wire \stat_rd_data_reg[9]_i_8_n_0 ;
  wire \stat_rd_data_reg[9]_i_9_n_0 ;
  wire [1:0]state;
  wire state15_out;
  wire state1__0;
  wire \state_reg_n_0_[0] ;
  wire \state_reg_n_0_[1] ;
  wire \tagged_frame_good[0]_i_2_n_0 ;
  wire [63:0]tagged_frame_good_reg;
  wire \tagged_frame_good_reg[0]_i_1_n_0 ;
  wire \tagged_frame_good_reg[0]_i_1_n_1 ;
  wire \tagged_frame_good_reg[0]_i_1_n_10 ;
  wire \tagged_frame_good_reg[0]_i_1_n_11 ;
  wire \tagged_frame_good_reg[0]_i_1_n_12 ;
  wire \tagged_frame_good_reg[0]_i_1_n_13 ;
  wire \tagged_frame_good_reg[0]_i_1_n_14 ;
  wire \tagged_frame_good_reg[0]_i_1_n_15 ;
  wire \tagged_frame_good_reg[0]_i_1_n_2 ;
  wire \tagged_frame_good_reg[0]_i_1_n_3 ;
  wire \tagged_frame_good_reg[0]_i_1_n_4 ;
  wire \tagged_frame_good_reg[0]_i_1_n_5 ;
  wire \tagged_frame_good_reg[0]_i_1_n_6 ;
  wire \tagged_frame_good_reg[0]_i_1_n_7 ;
  wire \tagged_frame_good_reg[0]_i_1_n_8 ;
  wire \tagged_frame_good_reg[0]_i_1_n_9 ;
  wire \tagged_frame_good_reg[16]_i_1_n_0 ;
  wire \tagged_frame_good_reg[16]_i_1_n_1 ;
  wire \tagged_frame_good_reg[16]_i_1_n_10 ;
  wire \tagged_frame_good_reg[16]_i_1_n_11 ;
  wire \tagged_frame_good_reg[16]_i_1_n_12 ;
  wire \tagged_frame_good_reg[16]_i_1_n_13 ;
  wire \tagged_frame_good_reg[16]_i_1_n_14 ;
  wire \tagged_frame_good_reg[16]_i_1_n_15 ;
  wire \tagged_frame_good_reg[16]_i_1_n_2 ;
  wire \tagged_frame_good_reg[16]_i_1_n_3 ;
  wire \tagged_frame_good_reg[16]_i_1_n_4 ;
  wire \tagged_frame_good_reg[16]_i_1_n_5 ;
  wire \tagged_frame_good_reg[16]_i_1_n_6 ;
  wire \tagged_frame_good_reg[16]_i_1_n_7 ;
  wire \tagged_frame_good_reg[16]_i_1_n_8 ;
  wire \tagged_frame_good_reg[16]_i_1_n_9 ;
  wire \tagged_frame_good_reg[24]_i_1_n_0 ;
  wire \tagged_frame_good_reg[24]_i_1_n_1 ;
  wire \tagged_frame_good_reg[24]_i_1_n_10 ;
  wire \tagged_frame_good_reg[24]_i_1_n_11 ;
  wire \tagged_frame_good_reg[24]_i_1_n_12 ;
  wire \tagged_frame_good_reg[24]_i_1_n_13 ;
  wire \tagged_frame_good_reg[24]_i_1_n_14 ;
  wire \tagged_frame_good_reg[24]_i_1_n_15 ;
  wire \tagged_frame_good_reg[24]_i_1_n_2 ;
  wire \tagged_frame_good_reg[24]_i_1_n_3 ;
  wire \tagged_frame_good_reg[24]_i_1_n_4 ;
  wire \tagged_frame_good_reg[24]_i_1_n_5 ;
  wire \tagged_frame_good_reg[24]_i_1_n_6 ;
  wire \tagged_frame_good_reg[24]_i_1_n_7 ;
  wire \tagged_frame_good_reg[24]_i_1_n_8 ;
  wire \tagged_frame_good_reg[24]_i_1_n_9 ;
  wire \tagged_frame_good_reg[32]_i_1_n_0 ;
  wire \tagged_frame_good_reg[32]_i_1_n_1 ;
  wire \tagged_frame_good_reg[32]_i_1_n_10 ;
  wire \tagged_frame_good_reg[32]_i_1_n_11 ;
  wire \tagged_frame_good_reg[32]_i_1_n_12 ;
  wire \tagged_frame_good_reg[32]_i_1_n_13 ;
  wire \tagged_frame_good_reg[32]_i_1_n_14 ;
  wire \tagged_frame_good_reg[32]_i_1_n_15 ;
  wire \tagged_frame_good_reg[32]_i_1_n_2 ;
  wire \tagged_frame_good_reg[32]_i_1_n_3 ;
  wire \tagged_frame_good_reg[32]_i_1_n_4 ;
  wire \tagged_frame_good_reg[32]_i_1_n_5 ;
  wire \tagged_frame_good_reg[32]_i_1_n_6 ;
  wire \tagged_frame_good_reg[32]_i_1_n_7 ;
  wire \tagged_frame_good_reg[32]_i_1_n_8 ;
  wire \tagged_frame_good_reg[32]_i_1_n_9 ;
  wire \tagged_frame_good_reg[40]_i_1_n_0 ;
  wire \tagged_frame_good_reg[40]_i_1_n_1 ;
  wire \tagged_frame_good_reg[40]_i_1_n_10 ;
  wire \tagged_frame_good_reg[40]_i_1_n_11 ;
  wire \tagged_frame_good_reg[40]_i_1_n_12 ;
  wire \tagged_frame_good_reg[40]_i_1_n_13 ;
  wire \tagged_frame_good_reg[40]_i_1_n_14 ;
  wire \tagged_frame_good_reg[40]_i_1_n_15 ;
  wire \tagged_frame_good_reg[40]_i_1_n_2 ;
  wire \tagged_frame_good_reg[40]_i_1_n_3 ;
  wire \tagged_frame_good_reg[40]_i_1_n_4 ;
  wire \tagged_frame_good_reg[40]_i_1_n_5 ;
  wire \tagged_frame_good_reg[40]_i_1_n_6 ;
  wire \tagged_frame_good_reg[40]_i_1_n_7 ;
  wire \tagged_frame_good_reg[40]_i_1_n_8 ;
  wire \tagged_frame_good_reg[40]_i_1_n_9 ;
  wire \tagged_frame_good_reg[48]_i_1_n_0 ;
  wire \tagged_frame_good_reg[48]_i_1_n_1 ;
  wire \tagged_frame_good_reg[48]_i_1_n_10 ;
  wire \tagged_frame_good_reg[48]_i_1_n_11 ;
  wire \tagged_frame_good_reg[48]_i_1_n_12 ;
  wire \tagged_frame_good_reg[48]_i_1_n_13 ;
  wire \tagged_frame_good_reg[48]_i_1_n_14 ;
  wire \tagged_frame_good_reg[48]_i_1_n_15 ;
  wire \tagged_frame_good_reg[48]_i_1_n_2 ;
  wire \tagged_frame_good_reg[48]_i_1_n_3 ;
  wire \tagged_frame_good_reg[48]_i_1_n_4 ;
  wire \tagged_frame_good_reg[48]_i_1_n_5 ;
  wire \tagged_frame_good_reg[48]_i_1_n_6 ;
  wire \tagged_frame_good_reg[48]_i_1_n_7 ;
  wire \tagged_frame_good_reg[48]_i_1_n_8 ;
  wire \tagged_frame_good_reg[48]_i_1_n_9 ;
  wire \tagged_frame_good_reg[56]_i_1_n_1 ;
  wire \tagged_frame_good_reg[56]_i_1_n_10 ;
  wire \tagged_frame_good_reg[56]_i_1_n_11 ;
  wire \tagged_frame_good_reg[56]_i_1_n_12 ;
  wire \tagged_frame_good_reg[56]_i_1_n_13 ;
  wire \tagged_frame_good_reg[56]_i_1_n_14 ;
  wire \tagged_frame_good_reg[56]_i_1_n_15 ;
  wire \tagged_frame_good_reg[56]_i_1_n_2 ;
  wire \tagged_frame_good_reg[56]_i_1_n_3 ;
  wire \tagged_frame_good_reg[56]_i_1_n_4 ;
  wire \tagged_frame_good_reg[56]_i_1_n_5 ;
  wire \tagged_frame_good_reg[56]_i_1_n_6 ;
  wire \tagged_frame_good_reg[56]_i_1_n_7 ;
  wire \tagged_frame_good_reg[56]_i_1_n_8 ;
  wire \tagged_frame_good_reg[56]_i_1_n_9 ;
  wire \tagged_frame_good_reg[8]_i_1_n_0 ;
  wire \tagged_frame_good_reg[8]_i_1_n_1 ;
  wire \tagged_frame_good_reg[8]_i_1_n_10 ;
  wire \tagged_frame_good_reg[8]_i_1_n_11 ;
  wire \tagged_frame_good_reg[8]_i_1_n_12 ;
  wire \tagged_frame_good_reg[8]_i_1_n_13 ;
  wire \tagged_frame_good_reg[8]_i_1_n_14 ;
  wire \tagged_frame_good_reg[8]_i_1_n_15 ;
  wire \tagged_frame_good_reg[8]_i_1_n_2 ;
  wire \tagged_frame_good_reg[8]_i_1_n_3 ;
  wire \tagged_frame_good_reg[8]_i_1_n_4 ;
  wire \tagged_frame_good_reg[8]_i_1_n_5 ;
  wire \tagged_frame_good_reg[8]_i_1_n_6 ;
  wire \tagged_frame_good_reg[8]_i_1_n_7 ;
  wire \tagged_frame_good_reg[8]_i_1_n_8 ;
  wire \tagged_frame_good_reg[8]_i_1_n_9 ;
  wire \tagged_frame_transed[0]_i_2_n_0 ;
  wire [63:0]tagged_frame_transed_reg;
  wire \tagged_frame_transed_reg[0]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[0]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[16]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[24]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[32]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[40]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[48]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[56]_i_1_n_9 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_0 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_1 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_10 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_11 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_12 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_13 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_14 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_15 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_2 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_3 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_4 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_5 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_6 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_7 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_8 ;
  wire \tagged_frame_transed_reg[8]_i_1_n_9 ;
  wire [4:0]tmp_cnt;
  wire \tmp_cnt[0]_i_1_n_0 ;
  wire \tmp_cnt[1]_i_1_n_0 ;
  wire \tmp_cnt[2]_i_1_n_0 ;
  wire \tmp_cnt[3]_i_1_n_0 ;
  wire \tmp_cnt[4]_i_1_n_0 ;
  wire \total_bytes_recved[0]_i_2_n_0 ;
  wire [63:0]total_bytes_recved_reg;
  wire \total_bytes_recved_reg[0]_i_1_n_0 ;
  wire \total_bytes_recved_reg[0]_i_1_n_1 ;
  wire \total_bytes_recved_reg[0]_i_1_n_10 ;
  wire \total_bytes_recved_reg[0]_i_1_n_11 ;
  wire \total_bytes_recved_reg[0]_i_1_n_12 ;
  wire \total_bytes_recved_reg[0]_i_1_n_13 ;
  wire \total_bytes_recved_reg[0]_i_1_n_14 ;
  wire \total_bytes_recved_reg[0]_i_1_n_15 ;
  wire \total_bytes_recved_reg[0]_i_1_n_2 ;
  wire \total_bytes_recved_reg[0]_i_1_n_3 ;
  wire \total_bytes_recved_reg[0]_i_1_n_4 ;
  wire \total_bytes_recved_reg[0]_i_1_n_5 ;
  wire \total_bytes_recved_reg[0]_i_1_n_6 ;
  wire \total_bytes_recved_reg[0]_i_1_n_7 ;
  wire \total_bytes_recved_reg[0]_i_1_n_8 ;
  wire \total_bytes_recved_reg[0]_i_1_n_9 ;
  wire \total_bytes_recved_reg[16]_i_1_n_0 ;
  wire \total_bytes_recved_reg[16]_i_1_n_1 ;
  wire \total_bytes_recved_reg[16]_i_1_n_10 ;
  wire \total_bytes_recved_reg[16]_i_1_n_11 ;
  wire \total_bytes_recved_reg[16]_i_1_n_12 ;
  wire \total_bytes_recved_reg[16]_i_1_n_13 ;
  wire \total_bytes_recved_reg[16]_i_1_n_14 ;
  wire \total_bytes_recved_reg[16]_i_1_n_15 ;
  wire \total_bytes_recved_reg[16]_i_1_n_2 ;
  wire \total_bytes_recved_reg[16]_i_1_n_3 ;
  wire \total_bytes_recved_reg[16]_i_1_n_4 ;
  wire \total_bytes_recved_reg[16]_i_1_n_5 ;
  wire \total_bytes_recved_reg[16]_i_1_n_6 ;
  wire \total_bytes_recved_reg[16]_i_1_n_7 ;
  wire \total_bytes_recved_reg[16]_i_1_n_8 ;
  wire \total_bytes_recved_reg[16]_i_1_n_9 ;
  wire \total_bytes_recved_reg[24]_i_1_n_0 ;
  wire \total_bytes_recved_reg[24]_i_1_n_1 ;
  wire \total_bytes_recved_reg[24]_i_1_n_10 ;
  wire \total_bytes_recved_reg[24]_i_1_n_11 ;
  wire \total_bytes_recved_reg[24]_i_1_n_12 ;
  wire \total_bytes_recved_reg[24]_i_1_n_13 ;
  wire \total_bytes_recved_reg[24]_i_1_n_14 ;
  wire \total_bytes_recved_reg[24]_i_1_n_15 ;
  wire \total_bytes_recved_reg[24]_i_1_n_2 ;
  wire \total_bytes_recved_reg[24]_i_1_n_3 ;
  wire \total_bytes_recved_reg[24]_i_1_n_4 ;
  wire \total_bytes_recved_reg[24]_i_1_n_5 ;
  wire \total_bytes_recved_reg[24]_i_1_n_6 ;
  wire \total_bytes_recved_reg[24]_i_1_n_7 ;
  wire \total_bytes_recved_reg[24]_i_1_n_8 ;
  wire \total_bytes_recved_reg[24]_i_1_n_9 ;
  wire \total_bytes_recved_reg[32]_i_1_n_0 ;
  wire \total_bytes_recved_reg[32]_i_1_n_1 ;
  wire \total_bytes_recved_reg[32]_i_1_n_10 ;
  wire \total_bytes_recved_reg[32]_i_1_n_11 ;
  wire \total_bytes_recved_reg[32]_i_1_n_12 ;
  wire \total_bytes_recved_reg[32]_i_1_n_13 ;
  wire \total_bytes_recved_reg[32]_i_1_n_14 ;
  wire \total_bytes_recved_reg[32]_i_1_n_15 ;
  wire \total_bytes_recved_reg[32]_i_1_n_2 ;
  wire \total_bytes_recved_reg[32]_i_1_n_3 ;
  wire \total_bytes_recved_reg[32]_i_1_n_4 ;
  wire \total_bytes_recved_reg[32]_i_1_n_5 ;
  wire \total_bytes_recved_reg[32]_i_1_n_6 ;
  wire \total_bytes_recved_reg[32]_i_1_n_7 ;
  wire \total_bytes_recved_reg[32]_i_1_n_8 ;
  wire \total_bytes_recved_reg[32]_i_1_n_9 ;
  wire \total_bytes_recved_reg[40]_i_1_n_0 ;
  wire \total_bytes_recved_reg[40]_i_1_n_1 ;
  wire \total_bytes_recved_reg[40]_i_1_n_10 ;
  wire \total_bytes_recved_reg[40]_i_1_n_11 ;
  wire \total_bytes_recved_reg[40]_i_1_n_12 ;
  wire \total_bytes_recved_reg[40]_i_1_n_13 ;
  wire \total_bytes_recved_reg[40]_i_1_n_14 ;
  wire \total_bytes_recved_reg[40]_i_1_n_15 ;
  wire \total_bytes_recved_reg[40]_i_1_n_2 ;
  wire \total_bytes_recved_reg[40]_i_1_n_3 ;
  wire \total_bytes_recved_reg[40]_i_1_n_4 ;
  wire \total_bytes_recved_reg[40]_i_1_n_5 ;
  wire \total_bytes_recved_reg[40]_i_1_n_6 ;
  wire \total_bytes_recved_reg[40]_i_1_n_7 ;
  wire \total_bytes_recved_reg[40]_i_1_n_8 ;
  wire \total_bytes_recved_reg[40]_i_1_n_9 ;
  wire \total_bytes_recved_reg[48]_i_1_n_0 ;
  wire \total_bytes_recved_reg[48]_i_1_n_1 ;
  wire \total_bytes_recved_reg[48]_i_1_n_10 ;
  wire \total_bytes_recved_reg[48]_i_1_n_11 ;
  wire \total_bytes_recved_reg[48]_i_1_n_12 ;
  wire \total_bytes_recved_reg[48]_i_1_n_13 ;
  wire \total_bytes_recved_reg[48]_i_1_n_14 ;
  wire \total_bytes_recved_reg[48]_i_1_n_15 ;
  wire \total_bytes_recved_reg[48]_i_1_n_2 ;
  wire \total_bytes_recved_reg[48]_i_1_n_3 ;
  wire \total_bytes_recved_reg[48]_i_1_n_4 ;
  wire \total_bytes_recved_reg[48]_i_1_n_5 ;
  wire \total_bytes_recved_reg[48]_i_1_n_6 ;
  wire \total_bytes_recved_reg[48]_i_1_n_7 ;
  wire \total_bytes_recved_reg[48]_i_1_n_8 ;
  wire \total_bytes_recved_reg[48]_i_1_n_9 ;
  wire \total_bytes_recved_reg[56]_i_1_n_1 ;
  wire \total_bytes_recved_reg[56]_i_1_n_10 ;
  wire \total_bytes_recved_reg[56]_i_1_n_11 ;
  wire \total_bytes_recved_reg[56]_i_1_n_12 ;
  wire \total_bytes_recved_reg[56]_i_1_n_13 ;
  wire \total_bytes_recved_reg[56]_i_1_n_14 ;
  wire \total_bytes_recved_reg[56]_i_1_n_15 ;
  wire \total_bytes_recved_reg[56]_i_1_n_2 ;
  wire \total_bytes_recved_reg[56]_i_1_n_3 ;
  wire \total_bytes_recved_reg[56]_i_1_n_4 ;
  wire \total_bytes_recved_reg[56]_i_1_n_5 ;
  wire \total_bytes_recved_reg[56]_i_1_n_6 ;
  wire \total_bytes_recved_reg[56]_i_1_n_7 ;
  wire \total_bytes_recved_reg[56]_i_1_n_8 ;
  wire \total_bytes_recved_reg[56]_i_1_n_9 ;
  wire \total_bytes_recved_reg[8]_i_1_n_0 ;
  wire \total_bytes_recved_reg[8]_i_1_n_1 ;
  wire \total_bytes_recved_reg[8]_i_1_n_10 ;
  wire \total_bytes_recved_reg[8]_i_1_n_11 ;
  wire \total_bytes_recved_reg[8]_i_1_n_12 ;
  wire \total_bytes_recved_reg[8]_i_1_n_13 ;
  wire \total_bytes_recved_reg[8]_i_1_n_14 ;
  wire \total_bytes_recved_reg[8]_i_1_n_15 ;
  wire \total_bytes_recved_reg[8]_i_1_n_2 ;
  wire \total_bytes_recved_reg[8]_i_1_n_3 ;
  wire \total_bytes_recved_reg[8]_i_1_n_4 ;
  wire \total_bytes_recved_reg[8]_i_1_n_5 ;
  wire \total_bytes_recved_reg[8]_i_1_n_6 ;
  wire \total_bytes_recved_reg[8]_i_1_n_7 ;
  wire \total_bytes_recved_reg[8]_i_1_n_8 ;
  wire \total_bytes_recved_reg[8]_i_1_n_9 ;
  wire \total_bytes_transed[0]_i_2_n_0 ;
  wire [63:0]total_bytes_transed_reg;
  wire \total_bytes_transed_reg[0]_i_1_n_0 ;
  wire \total_bytes_transed_reg[0]_i_1_n_1 ;
  wire \total_bytes_transed_reg[0]_i_1_n_10 ;
  wire \total_bytes_transed_reg[0]_i_1_n_11 ;
  wire \total_bytes_transed_reg[0]_i_1_n_12 ;
  wire \total_bytes_transed_reg[0]_i_1_n_13 ;
  wire \total_bytes_transed_reg[0]_i_1_n_14 ;
  wire \total_bytes_transed_reg[0]_i_1_n_15 ;
  wire \total_bytes_transed_reg[0]_i_1_n_2 ;
  wire \total_bytes_transed_reg[0]_i_1_n_3 ;
  wire \total_bytes_transed_reg[0]_i_1_n_4 ;
  wire \total_bytes_transed_reg[0]_i_1_n_5 ;
  wire \total_bytes_transed_reg[0]_i_1_n_6 ;
  wire \total_bytes_transed_reg[0]_i_1_n_7 ;
  wire \total_bytes_transed_reg[0]_i_1_n_8 ;
  wire \total_bytes_transed_reg[0]_i_1_n_9 ;
  wire \total_bytes_transed_reg[16]_i_1_n_0 ;
  wire \total_bytes_transed_reg[16]_i_1_n_1 ;
  wire \total_bytes_transed_reg[16]_i_1_n_10 ;
  wire \total_bytes_transed_reg[16]_i_1_n_11 ;
  wire \total_bytes_transed_reg[16]_i_1_n_12 ;
  wire \total_bytes_transed_reg[16]_i_1_n_13 ;
  wire \total_bytes_transed_reg[16]_i_1_n_14 ;
  wire \total_bytes_transed_reg[16]_i_1_n_15 ;
  wire \total_bytes_transed_reg[16]_i_1_n_2 ;
  wire \total_bytes_transed_reg[16]_i_1_n_3 ;
  wire \total_bytes_transed_reg[16]_i_1_n_4 ;
  wire \total_bytes_transed_reg[16]_i_1_n_5 ;
  wire \total_bytes_transed_reg[16]_i_1_n_6 ;
  wire \total_bytes_transed_reg[16]_i_1_n_7 ;
  wire \total_bytes_transed_reg[16]_i_1_n_8 ;
  wire \total_bytes_transed_reg[16]_i_1_n_9 ;
  wire \total_bytes_transed_reg[24]_i_1_n_0 ;
  wire \total_bytes_transed_reg[24]_i_1_n_1 ;
  wire \total_bytes_transed_reg[24]_i_1_n_10 ;
  wire \total_bytes_transed_reg[24]_i_1_n_11 ;
  wire \total_bytes_transed_reg[24]_i_1_n_12 ;
  wire \total_bytes_transed_reg[24]_i_1_n_13 ;
  wire \total_bytes_transed_reg[24]_i_1_n_14 ;
  wire \total_bytes_transed_reg[24]_i_1_n_15 ;
  wire \total_bytes_transed_reg[24]_i_1_n_2 ;
  wire \total_bytes_transed_reg[24]_i_1_n_3 ;
  wire \total_bytes_transed_reg[24]_i_1_n_4 ;
  wire \total_bytes_transed_reg[24]_i_1_n_5 ;
  wire \total_bytes_transed_reg[24]_i_1_n_6 ;
  wire \total_bytes_transed_reg[24]_i_1_n_7 ;
  wire \total_bytes_transed_reg[24]_i_1_n_8 ;
  wire \total_bytes_transed_reg[24]_i_1_n_9 ;
  wire \total_bytes_transed_reg[32]_i_1_n_0 ;
  wire \total_bytes_transed_reg[32]_i_1_n_1 ;
  wire \total_bytes_transed_reg[32]_i_1_n_10 ;
  wire \total_bytes_transed_reg[32]_i_1_n_11 ;
  wire \total_bytes_transed_reg[32]_i_1_n_12 ;
  wire \total_bytes_transed_reg[32]_i_1_n_13 ;
  wire \total_bytes_transed_reg[32]_i_1_n_14 ;
  wire \total_bytes_transed_reg[32]_i_1_n_15 ;
  wire \total_bytes_transed_reg[32]_i_1_n_2 ;
  wire \total_bytes_transed_reg[32]_i_1_n_3 ;
  wire \total_bytes_transed_reg[32]_i_1_n_4 ;
  wire \total_bytes_transed_reg[32]_i_1_n_5 ;
  wire \total_bytes_transed_reg[32]_i_1_n_6 ;
  wire \total_bytes_transed_reg[32]_i_1_n_7 ;
  wire \total_bytes_transed_reg[32]_i_1_n_8 ;
  wire \total_bytes_transed_reg[32]_i_1_n_9 ;
  wire \total_bytes_transed_reg[40]_i_1_n_0 ;
  wire \total_bytes_transed_reg[40]_i_1_n_1 ;
  wire \total_bytes_transed_reg[40]_i_1_n_10 ;
  wire \total_bytes_transed_reg[40]_i_1_n_11 ;
  wire \total_bytes_transed_reg[40]_i_1_n_12 ;
  wire \total_bytes_transed_reg[40]_i_1_n_13 ;
  wire \total_bytes_transed_reg[40]_i_1_n_14 ;
  wire \total_bytes_transed_reg[40]_i_1_n_15 ;
  wire \total_bytes_transed_reg[40]_i_1_n_2 ;
  wire \total_bytes_transed_reg[40]_i_1_n_3 ;
  wire \total_bytes_transed_reg[40]_i_1_n_4 ;
  wire \total_bytes_transed_reg[40]_i_1_n_5 ;
  wire \total_bytes_transed_reg[40]_i_1_n_6 ;
  wire \total_bytes_transed_reg[40]_i_1_n_7 ;
  wire \total_bytes_transed_reg[40]_i_1_n_8 ;
  wire \total_bytes_transed_reg[40]_i_1_n_9 ;
  wire \total_bytes_transed_reg[48]_i_1_n_0 ;
  wire \total_bytes_transed_reg[48]_i_1_n_1 ;
  wire \total_bytes_transed_reg[48]_i_1_n_10 ;
  wire \total_bytes_transed_reg[48]_i_1_n_11 ;
  wire \total_bytes_transed_reg[48]_i_1_n_12 ;
  wire \total_bytes_transed_reg[48]_i_1_n_13 ;
  wire \total_bytes_transed_reg[48]_i_1_n_14 ;
  wire \total_bytes_transed_reg[48]_i_1_n_15 ;
  wire \total_bytes_transed_reg[48]_i_1_n_2 ;
  wire \total_bytes_transed_reg[48]_i_1_n_3 ;
  wire \total_bytes_transed_reg[48]_i_1_n_4 ;
  wire \total_bytes_transed_reg[48]_i_1_n_5 ;
  wire \total_bytes_transed_reg[48]_i_1_n_6 ;
  wire \total_bytes_transed_reg[48]_i_1_n_7 ;
  wire \total_bytes_transed_reg[48]_i_1_n_8 ;
  wire \total_bytes_transed_reg[48]_i_1_n_9 ;
  wire \total_bytes_transed_reg[56]_i_1_n_1 ;
  wire \total_bytes_transed_reg[56]_i_1_n_10 ;
  wire \total_bytes_transed_reg[56]_i_1_n_11 ;
  wire \total_bytes_transed_reg[56]_i_1_n_12 ;
  wire \total_bytes_transed_reg[56]_i_1_n_13 ;
  wire \total_bytes_transed_reg[56]_i_1_n_14 ;
  wire \total_bytes_transed_reg[56]_i_1_n_15 ;
  wire \total_bytes_transed_reg[56]_i_1_n_2 ;
  wire \total_bytes_transed_reg[56]_i_1_n_3 ;
  wire \total_bytes_transed_reg[56]_i_1_n_4 ;
  wire \total_bytes_transed_reg[56]_i_1_n_5 ;
  wire \total_bytes_transed_reg[56]_i_1_n_6 ;
  wire \total_bytes_transed_reg[56]_i_1_n_7 ;
  wire \total_bytes_transed_reg[56]_i_1_n_8 ;
  wire \total_bytes_transed_reg[56]_i_1_n_9 ;
  wire \total_bytes_transed_reg[8]_i_1_n_0 ;
  wire \total_bytes_transed_reg[8]_i_1_n_1 ;
  wire \total_bytes_transed_reg[8]_i_1_n_10 ;
  wire \total_bytes_transed_reg[8]_i_1_n_11 ;
  wire \total_bytes_transed_reg[8]_i_1_n_12 ;
  wire \total_bytes_transed_reg[8]_i_1_n_13 ;
  wire \total_bytes_transed_reg[8]_i_1_n_14 ;
  wire \total_bytes_transed_reg[8]_i_1_n_15 ;
  wire \total_bytes_transed_reg[8]_i_1_n_2 ;
  wire \total_bytes_transed_reg[8]_i_1_n_3 ;
  wire \total_bytes_transed_reg[8]_i_1_n_4 ;
  wire \total_bytes_transed_reg[8]_i_1_n_5 ;
  wire \total_bytes_transed_reg[8]_i_1_n_6 ;
  wire \total_bytes_transed_reg[8]_i_1_n_7 ;
  wire \total_bytes_transed_reg[8]_i_1_n_8 ;
  wire \total_bytes_transed_reg[8]_i_1_n_9 ;
  wire \trans_config[31]_i_1_n_0 ;
  wire \trans_config[31]_i_2_n_0 ;
  wire \trans_config_reg_n_0_[0] ;
  wire \trans_config_reg_n_0_[10] ;
  wire \trans_config_reg_n_0_[11] ;
  wire \trans_config_reg_n_0_[12] ;
  wire \trans_config_reg_n_0_[13] ;
  wire \trans_config_reg_n_0_[14] ;
  wire \trans_config_reg_n_0_[15] ;
  wire \trans_config_reg_n_0_[16] ;
  wire \trans_config_reg_n_0_[17] ;
  wire \trans_config_reg_n_0_[18] ;
  wire \trans_config_reg_n_0_[19] ;
  wire \trans_config_reg_n_0_[1] ;
  wire \trans_config_reg_n_0_[20] ;
  wire \trans_config_reg_n_0_[21] ;
  wire \trans_config_reg_n_0_[22] ;
  wire \trans_config_reg_n_0_[23] ;
  wire \trans_config_reg_n_0_[2] ;
  wire \trans_config_reg_n_0_[3] ;
  wire \trans_config_reg_n_0_[4] ;
  wire \trans_config_reg_n_0_[5] ;
  wire \trans_config_reg_n_0_[6] ;
  wire \trans_config_reg_n_0_[7] ;
  wire \trans_config_reg_n_0_[8] ;
  wire \trans_config_reg_n_0_[9] ;
  wire [14:0]txStatRegPlus;
  wire \underrun_error[0]_i_2_n_0 ;
  wire [63:0]underrun_error_reg;
  wire \underrun_error_reg[0]_i_1_n_0 ;
  wire \underrun_error_reg[0]_i_1_n_1 ;
  wire \underrun_error_reg[0]_i_1_n_10 ;
  wire \underrun_error_reg[0]_i_1_n_11 ;
  wire \underrun_error_reg[0]_i_1_n_12 ;
  wire \underrun_error_reg[0]_i_1_n_13 ;
  wire \underrun_error_reg[0]_i_1_n_14 ;
  wire \underrun_error_reg[0]_i_1_n_15 ;
  wire \underrun_error_reg[0]_i_1_n_2 ;
  wire \underrun_error_reg[0]_i_1_n_3 ;
  wire \underrun_error_reg[0]_i_1_n_4 ;
  wire \underrun_error_reg[0]_i_1_n_5 ;
  wire \underrun_error_reg[0]_i_1_n_6 ;
  wire \underrun_error_reg[0]_i_1_n_7 ;
  wire \underrun_error_reg[0]_i_1_n_8 ;
  wire \underrun_error_reg[0]_i_1_n_9 ;
  wire \underrun_error_reg[16]_i_1_n_0 ;
  wire \underrun_error_reg[16]_i_1_n_1 ;
  wire \underrun_error_reg[16]_i_1_n_10 ;
  wire \underrun_error_reg[16]_i_1_n_11 ;
  wire \underrun_error_reg[16]_i_1_n_12 ;
  wire \underrun_error_reg[16]_i_1_n_13 ;
  wire \underrun_error_reg[16]_i_1_n_14 ;
  wire \underrun_error_reg[16]_i_1_n_15 ;
  wire \underrun_error_reg[16]_i_1_n_2 ;
  wire \underrun_error_reg[16]_i_1_n_3 ;
  wire \underrun_error_reg[16]_i_1_n_4 ;
  wire \underrun_error_reg[16]_i_1_n_5 ;
  wire \underrun_error_reg[16]_i_1_n_6 ;
  wire \underrun_error_reg[16]_i_1_n_7 ;
  wire \underrun_error_reg[16]_i_1_n_8 ;
  wire \underrun_error_reg[16]_i_1_n_9 ;
  wire \underrun_error_reg[24]_i_1_n_0 ;
  wire \underrun_error_reg[24]_i_1_n_1 ;
  wire \underrun_error_reg[24]_i_1_n_10 ;
  wire \underrun_error_reg[24]_i_1_n_11 ;
  wire \underrun_error_reg[24]_i_1_n_12 ;
  wire \underrun_error_reg[24]_i_1_n_13 ;
  wire \underrun_error_reg[24]_i_1_n_14 ;
  wire \underrun_error_reg[24]_i_1_n_15 ;
  wire \underrun_error_reg[24]_i_1_n_2 ;
  wire \underrun_error_reg[24]_i_1_n_3 ;
  wire \underrun_error_reg[24]_i_1_n_4 ;
  wire \underrun_error_reg[24]_i_1_n_5 ;
  wire \underrun_error_reg[24]_i_1_n_6 ;
  wire \underrun_error_reg[24]_i_1_n_7 ;
  wire \underrun_error_reg[24]_i_1_n_8 ;
  wire \underrun_error_reg[24]_i_1_n_9 ;
  wire \underrun_error_reg[32]_i_1_n_0 ;
  wire \underrun_error_reg[32]_i_1_n_1 ;
  wire \underrun_error_reg[32]_i_1_n_10 ;
  wire \underrun_error_reg[32]_i_1_n_11 ;
  wire \underrun_error_reg[32]_i_1_n_12 ;
  wire \underrun_error_reg[32]_i_1_n_13 ;
  wire \underrun_error_reg[32]_i_1_n_14 ;
  wire \underrun_error_reg[32]_i_1_n_15 ;
  wire \underrun_error_reg[32]_i_1_n_2 ;
  wire \underrun_error_reg[32]_i_1_n_3 ;
  wire \underrun_error_reg[32]_i_1_n_4 ;
  wire \underrun_error_reg[32]_i_1_n_5 ;
  wire \underrun_error_reg[32]_i_1_n_6 ;
  wire \underrun_error_reg[32]_i_1_n_7 ;
  wire \underrun_error_reg[32]_i_1_n_8 ;
  wire \underrun_error_reg[32]_i_1_n_9 ;
  wire \underrun_error_reg[40]_i_1_n_0 ;
  wire \underrun_error_reg[40]_i_1_n_1 ;
  wire \underrun_error_reg[40]_i_1_n_10 ;
  wire \underrun_error_reg[40]_i_1_n_11 ;
  wire \underrun_error_reg[40]_i_1_n_12 ;
  wire \underrun_error_reg[40]_i_1_n_13 ;
  wire \underrun_error_reg[40]_i_1_n_14 ;
  wire \underrun_error_reg[40]_i_1_n_15 ;
  wire \underrun_error_reg[40]_i_1_n_2 ;
  wire \underrun_error_reg[40]_i_1_n_3 ;
  wire \underrun_error_reg[40]_i_1_n_4 ;
  wire \underrun_error_reg[40]_i_1_n_5 ;
  wire \underrun_error_reg[40]_i_1_n_6 ;
  wire \underrun_error_reg[40]_i_1_n_7 ;
  wire \underrun_error_reg[40]_i_1_n_8 ;
  wire \underrun_error_reg[40]_i_1_n_9 ;
  wire \underrun_error_reg[48]_i_1_n_0 ;
  wire \underrun_error_reg[48]_i_1_n_1 ;
  wire \underrun_error_reg[48]_i_1_n_10 ;
  wire \underrun_error_reg[48]_i_1_n_11 ;
  wire \underrun_error_reg[48]_i_1_n_12 ;
  wire \underrun_error_reg[48]_i_1_n_13 ;
  wire \underrun_error_reg[48]_i_1_n_14 ;
  wire \underrun_error_reg[48]_i_1_n_15 ;
  wire \underrun_error_reg[48]_i_1_n_2 ;
  wire \underrun_error_reg[48]_i_1_n_3 ;
  wire \underrun_error_reg[48]_i_1_n_4 ;
  wire \underrun_error_reg[48]_i_1_n_5 ;
  wire \underrun_error_reg[48]_i_1_n_6 ;
  wire \underrun_error_reg[48]_i_1_n_7 ;
  wire \underrun_error_reg[48]_i_1_n_8 ;
  wire \underrun_error_reg[48]_i_1_n_9 ;
  wire \underrun_error_reg[56]_i_1_n_1 ;
  wire \underrun_error_reg[56]_i_1_n_10 ;
  wire \underrun_error_reg[56]_i_1_n_11 ;
  wire \underrun_error_reg[56]_i_1_n_12 ;
  wire \underrun_error_reg[56]_i_1_n_13 ;
  wire \underrun_error_reg[56]_i_1_n_14 ;
  wire \underrun_error_reg[56]_i_1_n_15 ;
  wire \underrun_error_reg[56]_i_1_n_2 ;
  wire \underrun_error_reg[56]_i_1_n_3 ;
  wire \underrun_error_reg[56]_i_1_n_4 ;
  wire \underrun_error_reg[56]_i_1_n_5 ;
  wire \underrun_error_reg[56]_i_1_n_6 ;
  wire \underrun_error_reg[56]_i_1_n_7 ;
  wire \underrun_error_reg[56]_i_1_n_8 ;
  wire \underrun_error_reg[56]_i_1_n_9 ;
  wire \underrun_error_reg[8]_i_1_n_0 ;
  wire \underrun_error_reg[8]_i_1_n_1 ;
  wire \underrun_error_reg[8]_i_1_n_10 ;
  wire \underrun_error_reg[8]_i_1_n_11 ;
  wire \underrun_error_reg[8]_i_1_n_12 ;
  wire \underrun_error_reg[8]_i_1_n_13 ;
  wire \underrun_error_reg[8]_i_1_n_14 ;
  wire \underrun_error_reg[8]_i_1_n_15 ;
  wire \underrun_error_reg[8]_i_1_n_2 ;
  wire \underrun_error_reg[8]_i_1_n_3 ;
  wire \underrun_error_reg[8]_i_1_n_4 ;
  wire \underrun_error_reg[8]_i_1_n_5 ;
  wire \underrun_error_reg[8]_i_1_n_6 ;
  wire \underrun_error_reg[8]_i_1_n_7 ;
  wire \underrun_error_reg[8]_i_1_n_8 ;
  wire \underrun_error_reg[8]_i_1_n_9 ;
  wire \undersize_frame[0]_i_2_n_0 ;
  wire [63:0]undersize_frame_reg;
  wire \undersize_frame_reg[0]_i_1_n_0 ;
  wire \undersize_frame_reg[0]_i_1_n_1 ;
  wire \undersize_frame_reg[0]_i_1_n_10 ;
  wire \undersize_frame_reg[0]_i_1_n_11 ;
  wire \undersize_frame_reg[0]_i_1_n_12 ;
  wire \undersize_frame_reg[0]_i_1_n_13 ;
  wire \undersize_frame_reg[0]_i_1_n_14 ;
  wire \undersize_frame_reg[0]_i_1_n_15 ;
  wire \undersize_frame_reg[0]_i_1_n_2 ;
  wire \undersize_frame_reg[0]_i_1_n_3 ;
  wire \undersize_frame_reg[0]_i_1_n_4 ;
  wire \undersize_frame_reg[0]_i_1_n_5 ;
  wire \undersize_frame_reg[0]_i_1_n_6 ;
  wire \undersize_frame_reg[0]_i_1_n_7 ;
  wire \undersize_frame_reg[0]_i_1_n_8 ;
  wire \undersize_frame_reg[0]_i_1_n_9 ;
  wire \undersize_frame_reg[16]_i_1_n_0 ;
  wire \undersize_frame_reg[16]_i_1_n_1 ;
  wire \undersize_frame_reg[16]_i_1_n_10 ;
  wire \undersize_frame_reg[16]_i_1_n_11 ;
  wire \undersize_frame_reg[16]_i_1_n_12 ;
  wire \undersize_frame_reg[16]_i_1_n_13 ;
  wire \undersize_frame_reg[16]_i_1_n_14 ;
  wire \undersize_frame_reg[16]_i_1_n_15 ;
  wire \undersize_frame_reg[16]_i_1_n_2 ;
  wire \undersize_frame_reg[16]_i_1_n_3 ;
  wire \undersize_frame_reg[16]_i_1_n_4 ;
  wire \undersize_frame_reg[16]_i_1_n_5 ;
  wire \undersize_frame_reg[16]_i_1_n_6 ;
  wire \undersize_frame_reg[16]_i_1_n_7 ;
  wire \undersize_frame_reg[16]_i_1_n_8 ;
  wire \undersize_frame_reg[16]_i_1_n_9 ;
  wire \undersize_frame_reg[24]_i_1_n_0 ;
  wire \undersize_frame_reg[24]_i_1_n_1 ;
  wire \undersize_frame_reg[24]_i_1_n_10 ;
  wire \undersize_frame_reg[24]_i_1_n_11 ;
  wire \undersize_frame_reg[24]_i_1_n_12 ;
  wire \undersize_frame_reg[24]_i_1_n_13 ;
  wire \undersize_frame_reg[24]_i_1_n_14 ;
  wire \undersize_frame_reg[24]_i_1_n_15 ;
  wire \undersize_frame_reg[24]_i_1_n_2 ;
  wire \undersize_frame_reg[24]_i_1_n_3 ;
  wire \undersize_frame_reg[24]_i_1_n_4 ;
  wire \undersize_frame_reg[24]_i_1_n_5 ;
  wire \undersize_frame_reg[24]_i_1_n_6 ;
  wire \undersize_frame_reg[24]_i_1_n_7 ;
  wire \undersize_frame_reg[24]_i_1_n_8 ;
  wire \undersize_frame_reg[24]_i_1_n_9 ;
  wire \undersize_frame_reg[32]_i_1_n_0 ;
  wire \undersize_frame_reg[32]_i_1_n_1 ;
  wire \undersize_frame_reg[32]_i_1_n_10 ;
  wire \undersize_frame_reg[32]_i_1_n_11 ;
  wire \undersize_frame_reg[32]_i_1_n_12 ;
  wire \undersize_frame_reg[32]_i_1_n_13 ;
  wire \undersize_frame_reg[32]_i_1_n_14 ;
  wire \undersize_frame_reg[32]_i_1_n_15 ;
  wire \undersize_frame_reg[32]_i_1_n_2 ;
  wire \undersize_frame_reg[32]_i_1_n_3 ;
  wire \undersize_frame_reg[32]_i_1_n_4 ;
  wire \undersize_frame_reg[32]_i_1_n_5 ;
  wire \undersize_frame_reg[32]_i_1_n_6 ;
  wire \undersize_frame_reg[32]_i_1_n_7 ;
  wire \undersize_frame_reg[32]_i_1_n_8 ;
  wire \undersize_frame_reg[32]_i_1_n_9 ;
  wire \undersize_frame_reg[40]_i_1_n_0 ;
  wire \undersize_frame_reg[40]_i_1_n_1 ;
  wire \undersize_frame_reg[40]_i_1_n_10 ;
  wire \undersize_frame_reg[40]_i_1_n_11 ;
  wire \undersize_frame_reg[40]_i_1_n_12 ;
  wire \undersize_frame_reg[40]_i_1_n_13 ;
  wire \undersize_frame_reg[40]_i_1_n_14 ;
  wire \undersize_frame_reg[40]_i_1_n_15 ;
  wire \undersize_frame_reg[40]_i_1_n_2 ;
  wire \undersize_frame_reg[40]_i_1_n_3 ;
  wire \undersize_frame_reg[40]_i_1_n_4 ;
  wire \undersize_frame_reg[40]_i_1_n_5 ;
  wire \undersize_frame_reg[40]_i_1_n_6 ;
  wire \undersize_frame_reg[40]_i_1_n_7 ;
  wire \undersize_frame_reg[40]_i_1_n_8 ;
  wire \undersize_frame_reg[40]_i_1_n_9 ;
  wire \undersize_frame_reg[48]_i_1_n_0 ;
  wire \undersize_frame_reg[48]_i_1_n_1 ;
  wire \undersize_frame_reg[48]_i_1_n_10 ;
  wire \undersize_frame_reg[48]_i_1_n_11 ;
  wire \undersize_frame_reg[48]_i_1_n_12 ;
  wire \undersize_frame_reg[48]_i_1_n_13 ;
  wire \undersize_frame_reg[48]_i_1_n_14 ;
  wire \undersize_frame_reg[48]_i_1_n_15 ;
  wire \undersize_frame_reg[48]_i_1_n_2 ;
  wire \undersize_frame_reg[48]_i_1_n_3 ;
  wire \undersize_frame_reg[48]_i_1_n_4 ;
  wire \undersize_frame_reg[48]_i_1_n_5 ;
  wire \undersize_frame_reg[48]_i_1_n_6 ;
  wire \undersize_frame_reg[48]_i_1_n_7 ;
  wire \undersize_frame_reg[48]_i_1_n_8 ;
  wire \undersize_frame_reg[48]_i_1_n_9 ;
  wire \undersize_frame_reg[56]_i_1_n_1 ;
  wire \undersize_frame_reg[56]_i_1_n_10 ;
  wire \undersize_frame_reg[56]_i_1_n_11 ;
  wire \undersize_frame_reg[56]_i_1_n_12 ;
  wire \undersize_frame_reg[56]_i_1_n_13 ;
  wire \undersize_frame_reg[56]_i_1_n_14 ;
  wire \undersize_frame_reg[56]_i_1_n_15 ;
  wire \undersize_frame_reg[56]_i_1_n_2 ;
  wire \undersize_frame_reg[56]_i_1_n_3 ;
  wire \undersize_frame_reg[56]_i_1_n_4 ;
  wire \undersize_frame_reg[56]_i_1_n_5 ;
  wire \undersize_frame_reg[56]_i_1_n_6 ;
  wire \undersize_frame_reg[56]_i_1_n_7 ;
  wire \undersize_frame_reg[56]_i_1_n_8 ;
  wire \undersize_frame_reg[56]_i_1_n_9 ;
  wire \undersize_frame_reg[8]_i_1_n_0 ;
  wire \undersize_frame_reg[8]_i_1_n_1 ;
  wire \undersize_frame_reg[8]_i_1_n_10 ;
  wire \undersize_frame_reg[8]_i_1_n_11 ;
  wire \undersize_frame_reg[8]_i_1_n_12 ;
  wire \undersize_frame_reg[8]_i_1_n_13 ;
  wire \undersize_frame_reg[8]_i_1_n_14 ;
  wire \undersize_frame_reg[8]_i_1_n_15 ;
  wire \undersize_frame_reg[8]_i_1_n_2 ;
  wire \undersize_frame_reg[8]_i_1_n_3 ;
  wire \undersize_frame_reg[8]_i_1_n_4 ;
  wire \undersize_frame_reg[8]_i_1_n_5 ;
  wire \undersize_frame_reg[8]_i_1_n_6 ;
  wire \undersize_frame_reg[8]_i_1_n_7 ;
  wire \undersize_frame_reg[8]_i_1_n_8 ;
  wire \undersize_frame_reg[8]_i_1_n_9 ;
  wire \unsupported_control_frame[0]_i_2_n_0 ;
  wire [63:0]unsupported_control_frame_reg;
  wire \unsupported_control_frame_reg[0]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[0]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[16]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[24]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[32]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[40]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[48]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[56]_i_1_n_9 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_0 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_1 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_10 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_11 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_12 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_13 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_14 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_15 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_2 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_3 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_4 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_5 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_6 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_7 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_8 ;
  wire \unsupported_control_frame_reg[8]_i_1_n_9 ;
  wire [7:7]\NLW_broadcast_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_broadcast_received_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_control_frame_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_control_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_fcs_error_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_fragment_frame_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_1024_max_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_1024_max_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_128_255_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_128_255_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_256_511_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_256_511_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_512_1023_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_512_1023_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_64_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_64_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_65_127_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_65_127_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_frame_received_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_good_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_lt_out_range_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_multicast_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_multicast_received_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_oversize_frame_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_oversize_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_pause_frame_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_pause_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_tagged_frame_good_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_tagged_frame_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_total_bytes_recved_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_total_bytes_transed_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_underrun_error_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_undersize_frame_reg[56]_i_1_CO_UNCONNECTED ;
  wire [7:7]\NLW_unsupported_control_frame_reg[56]_i_1_CO_UNCONNECTED ;

  LUT1 #(
    .INIT(2'h1)) 
    \broadcast_frame_transed[0]_i_2 
       (.I0(broadcast_frame_transed_reg[0]),
        .O(\broadcast_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[0]_i_1_n_0 ,\broadcast_frame_transed_reg[0]_i_1_n_1 ,\broadcast_frame_transed_reg[0]_i_1_n_2 ,\broadcast_frame_transed_reg[0]_i_1_n_3 ,\broadcast_frame_transed_reg[0]_i_1_n_4 ,\broadcast_frame_transed_reg[0]_i_1_n_5 ,\broadcast_frame_transed_reg[0]_i_1_n_6 ,\broadcast_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\broadcast_frame_transed_reg[0]_i_1_n_8 ,\broadcast_frame_transed_reg[0]_i_1_n_9 ,\broadcast_frame_transed_reg[0]_i_1_n_10 ,\broadcast_frame_transed_reg[0]_i_1_n_11 ,\broadcast_frame_transed_reg[0]_i_1_n_12 ,\broadcast_frame_transed_reg[0]_i_1_n_13 ,\broadcast_frame_transed_reg[0]_i_1_n_14 ,\broadcast_frame_transed_reg[0]_i_1_n_15 }),
        .S({broadcast_frame_transed_reg[7:1],\broadcast_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[16]_i_1 
       (.CI(\broadcast_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[16]_i_1_n_0 ,\broadcast_frame_transed_reg[16]_i_1_n_1 ,\broadcast_frame_transed_reg[16]_i_1_n_2 ,\broadcast_frame_transed_reg[16]_i_1_n_3 ,\broadcast_frame_transed_reg[16]_i_1_n_4 ,\broadcast_frame_transed_reg[16]_i_1_n_5 ,\broadcast_frame_transed_reg[16]_i_1_n_6 ,\broadcast_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[16]_i_1_n_8 ,\broadcast_frame_transed_reg[16]_i_1_n_9 ,\broadcast_frame_transed_reg[16]_i_1_n_10 ,\broadcast_frame_transed_reg[16]_i_1_n_11 ,\broadcast_frame_transed_reg[16]_i_1_n_12 ,\broadcast_frame_transed_reg[16]_i_1_n_13 ,\broadcast_frame_transed_reg[16]_i_1_n_14 ,\broadcast_frame_transed_reg[16]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[16]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[24]_i_1 
       (.CI(\broadcast_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[24]_i_1_n_0 ,\broadcast_frame_transed_reg[24]_i_1_n_1 ,\broadcast_frame_transed_reg[24]_i_1_n_2 ,\broadcast_frame_transed_reg[24]_i_1_n_3 ,\broadcast_frame_transed_reg[24]_i_1_n_4 ,\broadcast_frame_transed_reg[24]_i_1_n_5 ,\broadcast_frame_transed_reg[24]_i_1_n_6 ,\broadcast_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[24]_i_1_n_8 ,\broadcast_frame_transed_reg[24]_i_1_n_9 ,\broadcast_frame_transed_reg[24]_i_1_n_10 ,\broadcast_frame_transed_reg[24]_i_1_n_11 ,\broadcast_frame_transed_reg[24]_i_1_n_12 ,\broadcast_frame_transed_reg[24]_i_1_n_13 ,\broadcast_frame_transed_reg[24]_i_1_n_14 ,\broadcast_frame_transed_reg[24]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[24]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[32]_i_1 
       (.CI(\broadcast_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[32]_i_1_n_0 ,\broadcast_frame_transed_reg[32]_i_1_n_1 ,\broadcast_frame_transed_reg[32]_i_1_n_2 ,\broadcast_frame_transed_reg[32]_i_1_n_3 ,\broadcast_frame_transed_reg[32]_i_1_n_4 ,\broadcast_frame_transed_reg[32]_i_1_n_5 ,\broadcast_frame_transed_reg[32]_i_1_n_6 ,\broadcast_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[32]_i_1_n_8 ,\broadcast_frame_transed_reg[32]_i_1_n_9 ,\broadcast_frame_transed_reg[32]_i_1_n_10 ,\broadcast_frame_transed_reg[32]_i_1_n_11 ,\broadcast_frame_transed_reg[32]_i_1_n_12 ,\broadcast_frame_transed_reg[32]_i_1_n_13 ,\broadcast_frame_transed_reg[32]_i_1_n_14 ,\broadcast_frame_transed_reg[32]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[32]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[40]_i_1 
       (.CI(\broadcast_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[40]_i_1_n_0 ,\broadcast_frame_transed_reg[40]_i_1_n_1 ,\broadcast_frame_transed_reg[40]_i_1_n_2 ,\broadcast_frame_transed_reg[40]_i_1_n_3 ,\broadcast_frame_transed_reg[40]_i_1_n_4 ,\broadcast_frame_transed_reg[40]_i_1_n_5 ,\broadcast_frame_transed_reg[40]_i_1_n_6 ,\broadcast_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[40]_i_1_n_8 ,\broadcast_frame_transed_reg[40]_i_1_n_9 ,\broadcast_frame_transed_reg[40]_i_1_n_10 ,\broadcast_frame_transed_reg[40]_i_1_n_11 ,\broadcast_frame_transed_reg[40]_i_1_n_12 ,\broadcast_frame_transed_reg[40]_i_1_n_13 ,\broadcast_frame_transed_reg[40]_i_1_n_14 ,\broadcast_frame_transed_reg[40]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[40]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[48]_i_1 
       (.CI(\broadcast_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[48]_i_1_n_0 ,\broadcast_frame_transed_reg[48]_i_1_n_1 ,\broadcast_frame_transed_reg[48]_i_1_n_2 ,\broadcast_frame_transed_reg[48]_i_1_n_3 ,\broadcast_frame_transed_reg[48]_i_1_n_4 ,\broadcast_frame_transed_reg[48]_i_1_n_5 ,\broadcast_frame_transed_reg[48]_i_1_n_6 ,\broadcast_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[48]_i_1_n_8 ,\broadcast_frame_transed_reg[48]_i_1_n_9 ,\broadcast_frame_transed_reg[48]_i_1_n_10 ,\broadcast_frame_transed_reg[48]_i_1_n_11 ,\broadcast_frame_transed_reg[48]_i_1_n_12 ,\broadcast_frame_transed_reg[48]_i_1_n_13 ,\broadcast_frame_transed_reg[48]_i_1_n_14 ,\broadcast_frame_transed_reg[48]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[48]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[56]_i_1 
       (.CI(\broadcast_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_broadcast_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\broadcast_frame_transed_reg[56]_i_1_n_1 ,\broadcast_frame_transed_reg[56]_i_1_n_2 ,\broadcast_frame_transed_reg[56]_i_1_n_3 ,\broadcast_frame_transed_reg[56]_i_1_n_4 ,\broadcast_frame_transed_reg[56]_i_1_n_5 ,\broadcast_frame_transed_reg[56]_i_1_n_6 ,\broadcast_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[56]_i_1_n_8 ,\broadcast_frame_transed_reg[56]_i_1_n_9 ,\broadcast_frame_transed_reg[56]_i_1_n_10 ,\broadcast_frame_transed_reg[56]_i_1_n_11 ,\broadcast_frame_transed_reg[56]_i_1_n_12 ,\broadcast_frame_transed_reg[56]_i_1_n_13 ,\broadcast_frame_transed_reg[56]_i_1_n_14 ,\broadcast_frame_transed_reg[56]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_13 ),
        .Q(broadcast_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_12 ),
        .Q(broadcast_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_11 ),
        .Q(broadcast_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_10 ),
        .Q(broadcast_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[56]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_9 ),
        .Q(broadcast_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[0]_i_1_n_8 ),
        .Q(broadcast_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_15 ),
        .Q(broadcast_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_frame_transed_reg[8]_i_1 
       (.CI(\broadcast_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_frame_transed_reg[8]_i_1_n_0 ,\broadcast_frame_transed_reg[8]_i_1_n_1 ,\broadcast_frame_transed_reg[8]_i_1_n_2 ,\broadcast_frame_transed_reg[8]_i_1_n_3 ,\broadcast_frame_transed_reg[8]_i_1_n_4 ,\broadcast_frame_transed_reg[8]_i_1_n_5 ,\broadcast_frame_transed_reg[8]_i_1_n_6 ,\broadcast_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_frame_transed_reg[8]_i_1_n_8 ,\broadcast_frame_transed_reg[8]_i_1_n_9 ,\broadcast_frame_transed_reg[8]_i_1_n_10 ,\broadcast_frame_transed_reg[8]_i_1_n_11 ,\broadcast_frame_transed_reg[8]_i_1_n_12 ,\broadcast_frame_transed_reg[8]_i_1_n_13 ,\broadcast_frame_transed_reg[8]_i_1_n_14 ,\broadcast_frame_transed_reg[8]_i_1_n_15 }),
        .S(broadcast_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_frame_transed_reg[8]_i_1_n_14 ),
        .Q(broadcast_frame_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \broadcast_received_good[0]_i_2 
       (.I0(broadcast_received_good_reg[0]),
        .O(\broadcast_received_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[0]_i_1_n_0 ,\broadcast_received_good_reg[0]_i_1_n_1 ,\broadcast_received_good_reg[0]_i_1_n_2 ,\broadcast_received_good_reg[0]_i_1_n_3 ,\broadcast_received_good_reg[0]_i_1_n_4 ,\broadcast_received_good_reg[0]_i_1_n_5 ,\broadcast_received_good_reg[0]_i_1_n_6 ,\broadcast_received_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\broadcast_received_good_reg[0]_i_1_n_8 ,\broadcast_received_good_reg[0]_i_1_n_9 ,\broadcast_received_good_reg[0]_i_1_n_10 ,\broadcast_received_good_reg[0]_i_1_n_11 ,\broadcast_received_good_reg[0]_i_1_n_12 ,\broadcast_received_good_reg[0]_i_1_n_13 ,\broadcast_received_good_reg[0]_i_1_n_14 ,\broadcast_received_good_reg[0]_i_1_n_15 }),
        .S({broadcast_received_good_reg[7:1],\broadcast_received_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[16]_i_1 
       (.CI(\broadcast_received_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[16]_i_1_n_0 ,\broadcast_received_good_reg[16]_i_1_n_1 ,\broadcast_received_good_reg[16]_i_1_n_2 ,\broadcast_received_good_reg[16]_i_1_n_3 ,\broadcast_received_good_reg[16]_i_1_n_4 ,\broadcast_received_good_reg[16]_i_1_n_5 ,\broadcast_received_good_reg[16]_i_1_n_6 ,\broadcast_received_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[16]_i_1_n_8 ,\broadcast_received_good_reg[16]_i_1_n_9 ,\broadcast_received_good_reg[16]_i_1_n_10 ,\broadcast_received_good_reg[16]_i_1_n_11 ,\broadcast_received_good_reg[16]_i_1_n_12 ,\broadcast_received_good_reg[16]_i_1_n_13 ,\broadcast_received_good_reg[16]_i_1_n_14 ,\broadcast_received_good_reg[16]_i_1_n_15 }),
        .S(broadcast_received_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[16]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[24]_i_1 
       (.CI(\broadcast_received_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[24]_i_1_n_0 ,\broadcast_received_good_reg[24]_i_1_n_1 ,\broadcast_received_good_reg[24]_i_1_n_2 ,\broadcast_received_good_reg[24]_i_1_n_3 ,\broadcast_received_good_reg[24]_i_1_n_4 ,\broadcast_received_good_reg[24]_i_1_n_5 ,\broadcast_received_good_reg[24]_i_1_n_6 ,\broadcast_received_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[24]_i_1_n_8 ,\broadcast_received_good_reg[24]_i_1_n_9 ,\broadcast_received_good_reg[24]_i_1_n_10 ,\broadcast_received_good_reg[24]_i_1_n_11 ,\broadcast_received_good_reg[24]_i_1_n_12 ,\broadcast_received_good_reg[24]_i_1_n_13 ,\broadcast_received_good_reg[24]_i_1_n_14 ,\broadcast_received_good_reg[24]_i_1_n_15 }),
        .S(broadcast_received_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[24]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[32]_i_1 
       (.CI(\broadcast_received_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[32]_i_1_n_0 ,\broadcast_received_good_reg[32]_i_1_n_1 ,\broadcast_received_good_reg[32]_i_1_n_2 ,\broadcast_received_good_reg[32]_i_1_n_3 ,\broadcast_received_good_reg[32]_i_1_n_4 ,\broadcast_received_good_reg[32]_i_1_n_5 ,\broadcast_received_good_reg[32]_i_1_n_6 ,\broadcast_received_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[32]_i_1_n_8 ,\broadcast_received_good_reg[32]_i_1_n_9 ,\broadcast_received_good_reg[32]_i_1_n_10 ,\broadcast_received_good_reg[32]_i_1_n_11 ,\broadcast_received_good_reg[32]_i_1_n_12 ,\broadcast_received_good_reg[32]_i_1_n_13 ,\broadcast_received_good_reg[32]_i_1_n_14 ,\broadcast_received_good_reg[32]_i_1_n_15 }),
        .S(broadcast_received_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[32]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[40]_i_1 
       (.CI(\broadcast_received_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[40]_i_1_n_0 ,\broadcast_received_good_reg[40]_i_1_n_1 ,\broadcast_received_good_reg[40]_i_1_n_2 ,\broadcast_received_good_reg[40]_i_1_n_3 ,\broadcast_received_good_reg[40]_i_1_n_4 ,\broadcast_received_good_reg[40]_i_1_n_5 ,\broadcast_received_good_reg[40]_i_1_n_6 ,\broadcast_received_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[40]_i_1_n_8 ,\broadcast_received_good_reg[40]_i_1_n_9 ,\broadcast_received_good_reg[40]_i_1_n_10 ,\broadcast_received_good_reg[40]_i_1_n_11 ,\broadcast_received_good_reg[40]_i_1_n_12 ,\broadcast_received_good_reg[40]_i_1_n_13 ,\broadcast_received_good_reg[40]_i_1_n_14 ,\broadcast_received_good_reg[40]_i_1_n_15 }),
        .S(broadcast_received_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[40]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[48]_i_1 
       (.CI(\broadcast_received_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[48]_i_1_n_0 ,\broadcast_received_good_reg[48]_i_1_n_1 ,\broadcast_received_good_reg[48]_i_1_n_2 ,\broadcast_received_good_reg[48]_i_1_n_3 ,\broadcast_received_good_reg[48]_i_1_n_4 ,\broadcast_received_good_reg[48]_i_1_n_5 ,\broadcast_received_good_reg[48]_i_1_n_6 ,\broadcast_received_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[48]_i_1_n_8 ,\broadcast_received_good_reg[48]_i_1_n_9 ,\broadcast_received_good_reg[48]_i_1_n_10 ,\broadcast_received_good_reg[48]_i_1_n_11 ,\broadcast_received_good_reg[48]_i_1_n_12 ,\broadcast_received_good_reg[48]_i_1_n_13 ,\broadcast_received_good_reg[48]_i_1_n_14 ,\broadcast_received_good_reg[48]_i_1_n_15 }),
        .S(broadcast_received_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[48]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[56]_i_1 
       (.CI(\broadcast_received_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_broadcast_received_good_reg[56]_i_1_CO_UNCONNECTED [7],\broadcast_received_good_reg[56]_i_1_n_1 ,\broadcast_received_good_reg[56]_i_1_n_2 ,\broadcast_received_good_reg[56]_i_1_n_3 ,\broadcast_received_good_reg[56]_i_1_n_4 ,\broadcast_received_good_reg[56]_i_1_n_5 ,\broadcast_received_good_reg[56]_i_1_n_6 ,\broadcast_received_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[56]_i_1_n_8 ,\broadcast_received_good_reg[56]_i_1_n_9 ,\broadcast_received_good_reg[56]_i_1_n_10 ,\broadcast_received_good_reg[56]_i_1_n_11 ,\broadcast_received_good_reg[56]_i_1_n_12 ,\broadcast_received_good_reg[56]_i_1_n_13 ,\broadcast_received_good_reg[56]_i_1_n_14 ,\broadcast_received_good_reg[56]_i_1_n_15 }),
        .S(broadcast_received_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_13 ),
        .Q(broadcast_received_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_12 ),
        .Q(broadcast_received_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_11 ),
        .Q(broadcast_received_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_10 ),
        .Q(broadcast_received_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[56]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_9 ),
        .Q(broadcast_received_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[0]_i_1_n_8 ),
        .Q(broadcast_received_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_15 ),
        .Q(broadcast_received_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \broadcast_received_good_reg[8]_i_1 
       (.CI(\broadcast_received_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\broadcast_received_good_reg[8]_i_1_n_0 ,\broadcast_received_good_reg[8]_i_1_n_1 ,\broadcast_received_good_reg[8]_i_1_n_2 ,\broadcast_received_good_reg[8]_i_1_n_3 ,\broadcast_received_good_reg[8]_i_1_n_4 ,\broadcast_received_good_reg[8]_i_1_n_5 ,\broadcast_received_good_reg[8]_i_1_n_6 ,\broadcast_received_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\broadcast_received_good_reg[8]_i_1_n_8 ,\broadcast_received_good_reg[8]_i_1_n_9 ,\broadcast_received_good_reg[8]_i_1_n_10 ,\broadcast_received_good_reg[8]_i_1_n_11 ,\broadcast_received_good_reg[8]_i_1_n_12 ,\broadcast_received_good_reg[8]_i_1_n_13 ,\broadcast_received_good_reg[8]_i_1_n_14 ,\broadcast_received_good_reg[8]_i_1_n_15 }),
        .S(broadcast_received_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \broadcast_received_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[2]),
        .CLR(rst_i),
        .D(\broadcast_received_good_reg[8]_i_1_n_14 ),
        .Q(broadcast_received_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \control_frame_good[0]_i_2 
       (.I0(control_frame_good_reg[0]),
        .O(\control_frame_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_15 ),
        .Q(control_frame_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[0]_i_1_n_0 ,\control_frame_good_reg[0]_i_1_n_1 ,\control_frame_good_reg[0]_i_1_n_2 ,\control_frame_good_reg[0]_i_1_n_3 ,\control_frame_good_reg[0]_i_1_n_4 ,\control_frame_good_reg[0]_i_1_n_5 ,\control_frame_good_reg[0]_i_1_n_6 ,\control_frame_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\control_frame_good_reg[0]_i_1_n_8 ,\control_frame_good_reg[0]_i_1_n_9 ,\control_frame_good_reg[0]_i_1_n_10 ,\control_frame_good_reg[0]_i_1_n_11 ,\control_frame_good_reg[0]_i_1_n_12 ,\control_frame_good_reg[0]_i_1_n_13 ,\control_frame_good_reg[0]_i_1_n_14 ,\control_frame_good_reg[0]_i_1_n_15 }),
        .S({control_frame_good_reg[7:1],\control_frame_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_13 ),
        .Q(control_frame_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_12 ),
        .Q(control_frame_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_11 ),
        .Q(control_frame_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_10 ),
        .Q(control_frame_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_9 ),
        .Q(control_frame_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_8 ),
        .Q(control_frame_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_15 ),
        .Q(control_frame_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[16]_i_1 
       (.CI(\control_frame_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[16]_i_1_n_0 ,\control_frame_good_reg[16]_i_1_n_1 ,\control_frame_good_reg[16]_i_1_n_2 ,\control_frame_good_reg[16]_i_1_n_3 ,\control_frame_good_reg[16]_i_1_n_4 ,\control_frame_good_reg[16]_i_1_n_5 ,\control_frame_good_reg[16]_i_1_n_6 ,\control_frame_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[16]_i_1_n_8 ,\control_frame_good_reg[16]_i_1_n_9 ,\control_frame_good_reg[16]_i_1_n_10 ,\control_frame_good_reg[16]_i_1_n_11 ,\control_frame_good_reg[16]_i_1_n_12 ,\control_frame_good_reg[16]_i_1_n_13 ,\control_frame_good_reg[16]_i_1_n_14 ,\control_frame_good_reg[16]_i_1_n_15 }),
        .S(control_frame_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_14 ),
        .Q(control_frame_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_13 ),
        .Q(control_frame_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_12 ),
        .Q(control_frame_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_14 ),
        .Q(control_frame_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_11 ),
        .Q(control_frame_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_10 ),
        .Q(control_frame_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_9 ),
        .Q(control_frame_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[16]_i_1_n_8 ),
        .Q(control_frame_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_15 ),
        .Q(control_frame_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[24]_i_1 
       (.CI(\control_frame_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[24]_i_1_n_0 ,\control_frame_good_reg[24]_i_1_n_1 ,\control_frame_good_reg[24]_i_1_n_2 ,\control_frame_good_reg[24]_i_1_n_3 ,\control_frame_good_reg[24]_i_1_n_4 ,\control_frame_good_reg[24]_i_1_n_5 ,\control_frame_good_reg[24]_i_1_n_6 ,\control_frame_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[24]_i_1_n_8 ,\control_frame_good_reg[24]_i_1_n_9 ,\control_frame_good_reg[24]_i_1_n_10 ,\control_frame_good_reg[24]_i_1_n_11 ,\control_frame_good_reg[24]_i_1_n_12 ,\control_frame_good_reg[24]_i_1_n_13 ,\control_frame_good_reg[24]_i_1_n_14 ,\control_frame_good_reg[24]_i_1_n_15 }),
        .S(control_frame_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_14 ),
        .Q(control_frame_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_13 ),
        .Q(control_frame_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_12 ),
        .Q(control_frame_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_11 ),
        .Q(control_frame_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_10 ),
        .Q(control_frame_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_13 ),
        .Q(control_frame_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_9 ),
        .Q(control_frame_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[24]_i_1_n_8 ),
        .Q(control_frame_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_15 ),
        .Q(control_frame_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[32]_i_1 
       (.CI(\control_frame_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[32]_i_1_n_0 ,\control_frame_good_reg[32]_i_1_n_1 ,\control_frame_good_reg[32]_i_1_n_2 ,\control_frame_good_reg[32]_i_1_n_3 ,\control_frame_good_reg[32]_i_1_n_4 ,\control_frame_good_reg[32]_i_1_n_5 ,\control_frame_good_reg[32]_i_1_n_6 ,\control_frame_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[32]_i_1_n_8 ,\control_frame_good_reg[32]_i_1_n_9 ,\control_frame_good_reg[32]_i_1_n_10 ,\control_frame_good_reg[32]_i_1_n_11 ,\control_frame_good_reg[32]_i_1_n_12 ,\control_frame_good_reg[32]_i_1_n_13 ,\control_frame_good_reg[32]_i_1_n_14 ,\control_frame_good_reg[32]_i_1_n_15 }),
        .S(control_frame_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_14 ),
        .Q(control_frame_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_13 ),
        .Q(control_frame_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_12 ),
        .Q(control_frame_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_11 ),
        .Q(control_frame_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_10 ),
        .Q(control_frame_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_9 ),
        .Q(control_frame_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[32]_i_1_n_8 ),
        .Q(control_frame_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_12 ),
        .Q(control_frame_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_15 ),
        .Q(control_frame_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[40]_i_1 
       (.CI(\control_frame_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[40]_i_1_n_0 ,\control_frame_good_reg[40]_i_1_n_1 ,\control_frame_good_reg[40]_i_1_n_2 ,\control_frame_good_reg[40]_i_1_n_3 ,\control_frame_good_reg[40]_i_1_n_4 ,\control_frame_good_reg[40]_i_1_n_5 ,\control_frame_good_reg[40]_i_1_n_6 ,\control_frame_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[40]_i_1_n_8 ,\control_frame_good_reg[40]_i_1_n_9 ,\control_frame_good_reg[40]_i_1_n_10 ,\control_frame_good_reg[40]_i_1_n_11 ,\control_frame_good_reg[40]_i_1_n_12 ,\control_frame_good_reg[40]_i_1_n_13 ,\control_frame_good_reg[40]_i_1_n_14 ,\control_frame_good_reg[40]_i_1_n_15 }),
        .S(control_frame_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_14 ),
        .Q(control_frame_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_13 ),
        .Q(control_frame_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_12 ),
        .Q(control_frame_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_11 ),
        .Q(control_frame_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_10 ),
        .Q(control_frame_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_9 ),
        .Q(control_frame_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[40]_i_1_n_8 ),
        .Q(control_frame_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_15 ),
        .Q(control_frame_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[48]_i_1 
       (.CI(\control_frame_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[48]_i_1_n_0 ,\control_frame_good_reg[48]_i_1_n_1 ,\control_frame_good_reg[48]_i_1_n_2 ,\control_frame_good_reg[48]_i_1_n_3 ,\control_frame_good_reg[48]_i_1_n_4 ,\control_frame_good_reg[48]_i_1_n_5 ,\control_frame_good_reg[48]_i_1_n_6 ,\control_frame_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[48]_i_1_n_8 ,\control_frame_good_reg[48]_i_1_n_9 ,\control_frame_good_reg[48]_i_1_n_10 ,\control_frame_good_reg[48]_i_1_n_11 ,\control_frame_good_reg[48]_i_1_n_12 ,\control_frame_good_reg[48]_i_1_n_13 ,\control_frame_good_reg[48]_i_1_n_14 ,\control_frame_good_reg[48]_i_1_n_15 }),
        .S(control_frame_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_14 ),
        .Q(control_frame_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_11 ),
        .Q(control_frame_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_13 ),
        .Q(control_frame_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_12 ),
        .Q(control_frame_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_11 ),
        .Q(control_frame_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_10 ),
        .Q(control_frame_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_9 ),
        .Q(control_frame_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[48]_i_1_n_8 ),
        .Q(control_frame_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_15 ),
        .Q(control_frame_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[56]_i_1 
       (.CI(\control_frame_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_control_frame_good_reg[56]_i_1_CO_UNCONNECTED [7],\control_frame_good_reg[56]_i_1_n_1 ,\control_frame_good_reg[56]_i_1_n_2 ,\control_frame_good_reg[56]_i_1_n_3 ,\control_frame_good_reg[56]_i_1_n_4 ,\control_frame_good_reg[56]_i_1_n_5 ,\control_frame_good_reg[56]_i_1_n_6 ,\control_frame_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[56]_i_1_n_8 ,\control_frame_good_reg[56]_i_1_n_9 ,\control_frame_good_reg[56]_i_1_n_10 ,\control_frame_good_reg[56]_i_1_n_11 ,\control_frame_good_reg[56]_i_1_n_12 ,\control_frame_good_reg[56]_i_1_n_13 ,\control_frame_good_reg[56]_i_1_n_14 ,\control_frame_good_reg[56]_i_1_n_15 }),
        .S(control_frame_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_14 ),
        .Q(control_frame_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_13 ),
        .Q(control_frame_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_12 ),
        .Q(control_frame_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_10 ),
        .Q(control_frame_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_11 ),
        .Q(control_frame_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_10 ),
        .Q(control_frame_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_9 ),
        .Q(control_frame_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[56]_i_1_n_8 ),
        .Q(control_frame_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_9 ),
        .Q(control_frame_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[0]_i_1_n_8 ),
        .Q(control_frame_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_15 ),
        .Q(control_frame_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_good_reg[8]_i_1 
       (.CI(\control_frame_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_good_reg[8]_i_1_n_0 ,\control_frame_good_reg[8]_i_1_n_1 ,\control_frame_good_reg[8]_i_1_n_2 ,\control_frame_good_reg[8]_i_1_n_3 ,\control_frame_good_reg[8]_i_1_n_4 ,\control_frame_good_reg[8]_i_1_n_5 ,\control_frame_good_reg[8]_i_1_n_6 ,\control_frame_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_good_reg[8]_i_1_n_8 ,\control_frame_good_reg[8]_i_1_n_9 ,\control_frame_good_reg[8]_i_1_n_10 ,\control_frame_good_reg[8]_i_1_n_11 ,\control_frame_good_reg[8]_i_1_n_12 ,\control_frame_good_reg[8]_i_1_n_13 ,\control_frame_good_reg[8]_i_1_n_14 ,\control_frame_good_reg[8]_i_1_n_15 }),
        .S(control_frame_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[10]),
        .CLR(rst_i),
        .D(\control_frame_good_reg[8]_i_1_n_14 ),
        .Q(control_frame_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \control_frame_transed[0]_i_2 
       (.I0(control_frame_transed_reg[0]),
        .O(\control_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_15 ),
        .Q(control_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[0]_i_1_n_0 ,\control_frame_transed_reg[0]_i_1_n_1 ,\control_frame_transed_reg[0]_i_1_n_2 ,\control_frame_transed_reg[0]_i_1_n_3 ,\control_frame_transed_reg[0]_i_1_n_4 ,\control_frame_transed_reg[0]_i_1_n_5 ,\control_frame_transed_reg[0]_i_1_n_6 ,\control_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\control_frame_transed_reg[0]_i_1_n_8 ,\control_frame_transed_reg[0]_i_1_n_9 ,\control_frame_transed_reg[0]_i_1_n_10 ,\control_frame_transed_reg[0]_i_1_n_11 ,\control_frame_transed_reg[0]_i_1_n_12 ,\control_frame_transed_reg[0]_i_1_n_13 ,\control_frame_transed_reg[0]_i_1_n_14 ,\control_frame_transed_reg[0]_i_1_n_15 }),
        .S({control_frame_transed_reg[7:1],\control_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_13 ),
        .Q(control_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_12 ),
        .Q(control_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_11 ),
        .Q(control_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_10 ),
        .Q(control_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_9 ),
        .Q(control_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_8 ),
        .Q(control_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_15 ),
        .Q(control_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[16]_i_1 
       (.CI(\control_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[16]_i_1_n_0 ,\control_frame_transed_reg[16]_i_1_n_1 ,\control_frame_transed_reg[16]_i_1_n_2 ,\control_frame_transed_reg[16]_i_1_n_3 ,\control_frame_transed_reg[16]_i_1_n_4 ,\control_frame_transed_reg[16]_i_1_n_5 ,\control_frame_transed_reg[16]_i_1_n_6 ,\control_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[16]_i_1_n_8 ,\control_frame_transed_reg[16]_i_1_n_9 ,\control_frame_transed_reg[16]_i_1_n_10 ,\control_frame_transed_reg[16]_i_1_n_11 ,\control_frame_transed_reg[16]_i_1_n_12 ,\control_frame_transed_reg[16]_i_1_n_13 ,\control_frame_transed_reg[16]_i_1_n_14 ,\control_frame_transed_reg[16]_i_1_n_15 }),
        .S(control_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_14 ),
        .Q(control_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_13 ),
        .Q(control_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_12 ),
        .Q(control_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_14 ),
        .Q(control_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_11 ),
        .Q(control_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_10 ),
        .Q(control_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_9 ),
        .Q(control_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[16]_i_1_n_8 ),
        .Q(control_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_15 ),
        .Q(control_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[24]_i_1 
       (.CI(\control_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[24]_i_1_n_0 ,\control_frame_transed_reg[24]_i_1_n_1 ,\control_frame_transed_reg[24]_i_1_n_2 ,\control_frame_transed_reg[24]_i_1_n_3 ,\control_frame_transed_reg[24]_i_1_n_4 ,\control_frame_transed_reg[24]_i_1_n_5 ,\control_frame_transed_reg[24]_i_1_n_6 ,\control_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[24]_i_1_n_8 ,\control_frame_transed_reg[24]_i_1_n_9 ,\control_frame_transed_reg[24]_i_1_n_10 ,\control_frame_transed_reg[24]_i_1_n_11 ,\control_frame_transed_reg[24]_i_1_n_12 ,\control_frame_transed_reg[24]_i_1_n_13 ,\control_frame_transed_reg[24]_i_1_n_14 ,\control_frame_transed_reg[24]_i_1_n_15 }),
        .S(control_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_14 ),
        .Q(control_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_13 ),
        .Q(control_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_12 ),
        .Q(control_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_11 ),
        .Q(control_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_10 ),
        .Q(control_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_13 ),
        .Q(control_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_9 ),
        .Q(control_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[24]_i_1_n_8 ),
        .Q(control_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_15 ),
        .Q(control_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[32]_i_1 
       (.CI(\control_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[32]_i_1_n_0 ,\control_frame_transed_reg[32]_i_1_n_1 ,\control_frame_transed_reg[32]_i_1_n_2 ,\control_frame_transed_reg[32]_i_1_n_3 ,\control_frame_transed_reg[32]_i_1_n_4 ,\control_frame_transed_reg[32]_i_1_n_5 ,\control_frame_transed_reg[32]_i_1_n_6 ,\control_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[32]_i_1_n_8 ,\control_frame_transed_reg[32]_i_1_n_9 ,\control_frame_transed_reg[32]_i_1_n_10 ,\control_frame_transed_reg[32]_i_1_n_11 ,\control_frame_transed_reg[32]_i_1_n_12 ,\control_frame_transed_reg[32]_i_1_n_13 ,\control_frame_transed_reg[32]_i_1_n_14 ,\control_frame_transed_reg[32]_i_1_n_15 }),
        .S(control_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_14 ),
        .Q(control_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_13 ),
        .Q(control_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_12 ),
        .Q(control_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_11 ),
        .Q(control_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_10 ),
        .Q(control_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_9 ),
        .Q(control_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[32]_i_1_n_8 ),
        .Q(control_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_12 ),
        .Q(control_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_15 ),
        .Q(control_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[40]_i_1 
       (.CI(\control_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[40]_i_1_n_0 ,\control_frame_transed_reg[40]_i_1_n_1 ,\control_frame_transed_reg[40]_i_1_n_2 ,\control_frame_transed_reg[40]_i_1_n_3 ,\control_frame_transed_reg[40]_i_1_n_4 ,\control_frame_transed_reg[40]_i_1_n_5 ,\control_frame_transed_reg[40]_i_1_n_6 ,\control_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[40]_i_1_n_8 ,\control_frame_transed_reg[40]_i_1_n_9 ,\control_frame_transed_reg[40]_i_1_n_10 ,\control_frame_transed_reg[40]_i_1_n_11 ,\control_frame_transed_reg[40]_i_1_n_12 ,\control_frame_transed_reg[40]_i_1_n_13 ,\control_frame_transed_reg[40]_i_1_n_14 ,\control_frame_transed_reg[40]_i_1_n_15 }),
        .S(control_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_14 ),
        .Q(control_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_13 ),
        .Q(control_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_12 ),
        .Q(control_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_11 ),
        .Q(control_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_10 ),
        .Q(control_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_9 ),
        .Q(control_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[40]_i_1_n_8 ),
        .Q(control_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_15 ),
        .Q(control_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[48]_i_1 
       (.CI(\control_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[48]_i_1_n_0 ,\control_frame_transed_reg[48]_i_1_n_1 ,\control_frame_transed_reg[48]_i_1_n_2 ,\control_frame_transed_reg[48]_i_1_n_3 ,\control_frame_transed_reg[48]_i_1_n_4 ,\control_frame_transed_reg[48]_i_1_n_5 ,\control_frame_transed_reg[48]_i_1_n_6 ,\control_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[48]_i_1_n_8 ,\control_frame_transed_reg[48]_i_1_n_9 ,\control_frame_transed_reg[48]_i_1_n_10 ,\control_frame_transed_reg[48]_i_1_n_11 ,\control_frame_transed_reg[48]_i_1_n_12 ,\control_frame_transed_reg[48]_i_1_n_13 ,\control_frame_transed_reg[48]_i_1_n_14 ,\control_frame_transed_reg[48]_i_1_n_15 }),
        .S(control_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_14 ),
        .Q(control_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_11 ),
        .Q(control_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_13 ),
        .Q(control_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_12 ),
        .Q(control_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_11 ),
        .Q(control_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_10 ),
        .Q(control_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_9 ),
        .Q(control_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[48]_i_1_n_8 ),
        .Q(control_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_15 ),
        .Q(control_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[56]_i_1 
       (.CI(\control_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_control_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\control_frame_transed_reg[56]_i_1_n_1 ,\control_frame_transed_reg[56]_i_1_n_2 ,\control_frame_transed_reg[56]_i_1_n_3 ,\control_frame_transed_reg[56]_i_1_n_4 ,\control_frame_transed_reg[56]_i_1_n_5 ,\control_frame_transed_reg[56]_i_1_n_6 ,\control_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[56]_i_1_n_8 ,\control_frame_transed_reg[56]_i_1_n_9 ,\control_frame_transed_reg[56]_i_1_n_10 ,\control_frame_transed_reg[56]_i_1_n_11 ,\control_frame_transed_reg[56]_i_1_n_12 ,\control_frame_transed_reg[56]_i_1_n_13 ,\control_frame_transed_reg[56]_i_1_n_14 ,\control_frame_transed_reg[56]_i_1_n_15 }),
        .S(control_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_14 ),
        .Q(control_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_13 ),
        .Q(control_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_12 ),
        .Q(control_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_10 ),
        .Q(control_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_11 ),
        .Q(control_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_10 ),
        .Q(control_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_9 ),
        .Q(control_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[56]_i_1_n_8 ),
        .Q(control_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_9 ),
        .Q(control_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[0]_i_1_n_8 ),
        .Q(control_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_15 ),
        .Q(control_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \control_frame_transed_reg[8]_i_1 
       (.CI(\control_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\control_frame_transed_reg[8]_i_1_n_0 ,\control_frame_transed_reg[8]_i_1_n_1 ,\control_frame_transed_reg[8]_i_1_n_2 ,\control_frame_transed_reg[8]_i_1_n_3 ,\control_frame_transed_reg[8]_i_1_n_4 ,\control_frame_transed_reg[8]_i_1_n_5 ,\control_frame_transed_reg[8]_i_1_n_6 ,\control_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\control_frame_transed_reg[8]_i_1_n_8 ,\control_frame_transed_reg[8]_i_1_n_9 ,\control_frame_transed_reg[8]_i_1_n_10 ,\control_frame_transed_reg[8]_i_1_n_11 ,\control_frame_transed_reg[8]_i_1_n_12 ,\control_frame_transed_reg[8]_i_1_n_13 ,\control_frame_transed_reg[8]_i_1_n_14 ,\control_frame_transed_reg[8]_i_1_n_15 }),
        .S(control_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \control_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[5]),
        .CLR(rst_i),
        .D(\control_frame_transed_reg[8]_i_1_n_14 ),
        .Q(control_frame_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    data_sel_i_1
       (.I0(\state_reg_n_0_[0] ),
        .O(read_done));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT2 #(
    .INIT(4'h2)) 
    data_sel_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(data_sel),
        .O(data_sel_i_2_n_0));
  FDCE #(
    .INIT(1'b0)) 
    data_sel_reg
       (.C(clk_i),
        .CE(read_done),
        .CLR(rst_i),
        .D(data_sel_i_2_n_0),
        .Q(data_sel));
  LUT1 #(
    .INIT(2'h1)) 
    \fcs_error[0]_i_2 
       (.I0(fcs_error_reg[0]),
        .O(\fcs_error[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_15 ),
        .Q(fcs_error_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[0]_i_1_n_0 ,\fcs_error_reg[0]_i_1_n_1 ,\fcs_error_reg[0]_i_1_n_2 ,\fcs_error_reg[0]_i_1_n_3 ,\fcs_error_reg[0]_i_1_n_4 ,\fcs_error_reg[0]_i_1_n_5 ,\fcs_error_reg[0]_i_1_n_6 ,\fcs_error_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\fcs_error_reg[0]_i_1_n_8 ,\fcs_error_reg[0]_i_1_n_9 ,\fcs_error_reg[0]_i_1_n_10 ,\fcs_error_reg[0]_i_1_n_11 ,\fcs_error_reg[0]_i_1_n_12 ,\fcs_error_reg[0]_i_1_n_13 ,\fcs_error_reg[0]_i_1_n_14 ,\fcs_error_reg[0]_i_1_n_15 }),
        .S({fcs_error_reg[7:1],\fcs_error[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_13 ),
        .Q(fcs_error_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_12 ),
        .Q(fcs_error_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_11 ),
        .Q(fcs_error_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_10 ),
        .Q(fcs_error_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_9 ),
        .Q(fcs_error_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_8 ),
        .Q(fcs_error_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_15 ),
        .Q(fcs_error_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[16]_i_1 
       (.CI(\fcs_error_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[16]_i_1_n_0 ,\fcs_error_reg[16]_i_1_n_1 ,\fcs_error_reg[16]_i_1_n_2 ,\fcs_error_reg[16]_i_1_n_3 ,\fcs_error_reg[16]_i_1_n_4 ,\fcs_error_reg[16]_i_1_n_5 ,\fcs_error_reg[16]_i_1_n_6 ,\fcs_error_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[16]_i_1_n_8 ,\fcs_error_reg[16]_i_1_n_9 ,\fcs_error_reg[16]_i_1_n_10 ,\fcs_error_reg[16]_i_1_n_11 ,\fcs_error_reg[16]_i_1_n_12 ,\fcs_error_reg[16]_i_1_n_13 ,\fcs_error_reg[16]_i_1_n_14 ,\fcs_error_reg[16]_i_1_n_15 }),
        .S(fcs_error_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_14 ),
        .Q(fcs_error_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_13 ),
        .Q(fcs_error_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_12 ),
        .Q(fcs_error_reg[19]));
  FDPE #(
    .INIT(1'b1)) 
    \fcs_error_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .D(\fcs_error_reg[0]_i_1_n_14 ),
        .PRE(rst_i),
        .Q(fcs_error_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_11 ),
        .Q(fcs_error_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_10 ),
        .Q(fcs_error_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_9 ),
        .Q(fcs_error_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[16]_i_1_n_8 ),
        .Q(fcs_error_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_15 ),
        .Q(fcs_error_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[24]_i_1 
       (.CI(\fcs_error_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[24]_i_1_n_0 ,\fcs_error_reg[24]_i_1_n_1 ,\fcs_error_reg[24]_i_1_n_2 ,\fcs_error_reg[24]_i_1_n_3 ,\fcs_error_reg[24]_i_1_n_4 ,\fcs_error_reg[24]_i_1_n_5 ,\fcs_error_reg[24]_i_1_n_6 ,\fcs_error_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[24]_i_1_n_8 ,\fcs_error_reg[24]_i_1_n_9 ,\fcs_error_reg[24]_i_1_n_10 ,\fcs_error_reg[24]_i_1_n_11 ,\fcs_error_reg[24]_i_1_n_12 ,\fcs_error_reg[24]_i_1_n_13 ,\fcs_error_reg[24]_i_1_n_14 ,\fcs_error_reg[24]_i_1_n_15 }),
        .S(fcs_error_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_14 ),
        .Q(fcs_error_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_13 ),
        .Q(fcs_error_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_12 ),
        .Q(fcs_error_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_11 ),
        .Q(fcs_error_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_10 ),
        .Q(fcs_error_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_13 ),
        .Q(fcs_error_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_9 ),
        .Q(fcs_error_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[24]_i_1_n_8 ),
        .Q(fcs_error_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_15 ),
        .Q(fcs_error_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[32]_i_1 
       (.CI(\fcs_error_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[32]_i_1_n_0 ,\fcs_error_reg[32]_i_1_n_1 ,\fcs_error_reg[32]_i_1_n_2 ,\fcs_error_reg[32]_i_1_n_3 ,\fcs_error_reg[32]_i_1_n_4 ,\fcs_error_reg[32]_i_1_n_5 ,\fcs_error_reg[32]_i_1_n_6 ,\fcs_error_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[32]_i_1_n_8 ,\fcs_error_reg[32]_i_1_n_9 ,\fcs_error_reg[32]_i_1_n_10 ,\fcs_error_reg[32]_i_1_n_11 ,\fcs_error_reg[32]_i_1_n_12 ,\fcs_error_reg[32]_i_1_n_13 ,\fcs_error_reg[32]_i_1_n_14 ,\fcs_error_reg[32]_i_1_n_15 }),
        .S(fcs_error_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_14 ),
        .Q(fcs_error_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_13 ),
        .Q(fcs_error_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_12 ),
        .Q(fcs_error_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_11 ),
        .Q(fcs_error_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_10 ),
        .Q(fcs_error_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_9 ),
        .Q(fcs_error_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[32]_i_1_n_8 ),
        .Q(fcs_error_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_12 ),
        .Q(fcs_error_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_15 ),
        .Q(fcs_error_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[40]_i_1 
       (.CI(\fcs_error_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[40]_i_1_n_0 ,\fcs_error_reg[40]_i_1_n_1 ,\fcs_error_reg[40]_i_1_n_2 ,\fcs_error_reg[40]_i_1_n_3 ,\fcs_error_reg[40]_i_1_n_4 ,\fcs_error_reg[40]_i_1_n_5 ,\fcs_error_reg[40]_i_1_n_6 ,\fcs_error_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[40]_i_1_n_8 ,\fcs_error_reg[40]_i_1_n_9 ,\fcs_error_reg[40]_i_1_n_10 ,\fcs_error_reg[40]_i_1_n_11 ,\fcs_error_reg[40]_i_1_n_12 ,\fcs_error_reg[40]_i_1_n_13 ,\fcs_error_reg[40]_i_1_n_14 ,\fcs_error_reg[40]_i_1_n_15 }),
        .S(fcs_error_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_14 ),
        .Q(fcs_error_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_13 ),
        .Q(fcs_error_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_12 ),
        .Q(fcs_error_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_11 ),
        .Q(fcs_error_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_10 ),
        .Q(fcs_error_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_9 ),
        .Q(fcs_error_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[40]_i_1_n_8 ),
        .Q(fcs_error_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_15 ),
        .Q(fcs_error_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[48]_i_1 
       (.CI(\fcs_error_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[48]_i_1_n_0 ,\fcs_error_reg[48]_i_1_n_1 ,\fcs_error_reg[48]_i_1_n_2 ,\fcs_error_reg[48]_i_1_n_3 ,\fcs_error_reg[48]_i_1_n_4 ,\fcs_error_reg[48]_i_1_n_5 ,\fcs_error_reg[48]_i_1_n_6 ,\fcs_error_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[48]_i_1_n_8 ,\fcs_error_reg[48]_i_1_n_9 ,\fcs_error_reg[48]_i_1_n_10 ,\fcs_error_reg[48]_i_1_n_11 ,\fcs_error_reg[48]_i_1_n_12 ,\fcs_error_reg[48]_i_1_n_13 ,\fcs_error_reg[48]_i_1_n_14 ,\fcs_error_reg[48]_i_1_n_15 }),
        .S(fcs_error_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_14 ),
        .Q(fcs_error_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_11 ),
        .Q(fcs_error_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_13 ),
        .Q(fcs_error_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_12 ),
        .Q(fcs_error_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_11 ),
        .Q(fcs_error_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_10 ),
        .Q(fcs_error_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_9 ),
        .Q(fcs_error_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[48]_i_1_n_8 ),
        .Q(fcs_error_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_15 ),
        .Q(fcs_error_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[56]_i_1 
       (.CI(\fcs_error_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_fcs_error_reg[56]_i_1_CO_UNCONNECTED [7],\fcs_error_reg[56]_i_1_n_1 ,\fcs_error_reg[56]_i_1_n_2 ,\fcs_error_reg[56]_i_1_n_3 ,\fcs_error_reg[56]_i_1_n_4 ,\fcs_error_reg[56]_i_1_n_5 ,\fcs_error_reg[56]_i_1_n_6 ,\fcs_error_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[56]_i_1_n_8 ,\fcs_error_reg[56]_i_1_n_9 ,\fcs_error_reg[56]_i_1_n_10 ,\fcs_error_reg[56]_i_1_n_11 ,\fcs_error_reg[56]_i_1_n_12 ,\fcs_error_reg[56]_i_1_n_13 ,\fcs_error_reg[56]_i_1_n_14 ,\fcs_error_reg[56]_i_1_n_15 }),
        .S(fcs_error_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_14 ),
        .Q(fcs_error_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_13 ),
        .Q(fcs_error_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_12 ),
        .Q(fcs_error_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_10 ),
        .Q(fcs_error_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_11 ),
        .Q(fcs_error_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_10 ),
        .Q(fcs_error_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_9 ),
        .Q(fcs_error_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[56]_i_1_n_8 ),
        .Q(fcs_error_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_9 ),
        .Q(fcs_error_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[0]_i_1_n_8 ),
        .Q(fcs_error_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_15 ),
        .Q(fcs_error_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fcs_error_reg[8]_i_1 
       (.CI(\fcs_error_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fcs_error_reg[8]_i_1_n_0 ,\fcs_error_reg[8]_i_1_n_1 ,\fcs_error_reg[8]_i_1_n_2 ,\fcs_error_reg[8]_i_1_n_3 ,\fcs_error_reg[8]_i_1_n_4 ,\fcs_error_reg[8]_i_1_n_5 ,\fcs_error_reg[8]_i_1_n_6 ,\fcs_error_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fcs_error_reg[8]_i_1_n_8 ,\fcs_error_reg[8]_i_1_n_9 ,\fcs_error_reg[8]_i_1_n_10 ,\fcs_error_reg[8]_i_1_n_11 ,\fcs_error_reg[8]_i_1_n_12 ,\fcs_error_reg[8]_i_1_n_13 ,\fcs_error_reg[8]_i_1_n_14 ,\fcs_error_reg[8]_i_1_n_15 }),
        .S(fcs_error_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \fcs_error_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[1]),
        .CLR(rst_i),
        .D(\fcs_error_reg[8]_i_1_n_14 ),
        .Q(fcs_error_reg[9]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \flow_control_config[31]_i_1 
       (.I0(recv_config01__0),
        .I1(\recv_config1[31]_i_3_n_0 ),
        .I2(out[1]),
        .I3(out[8]),
        .I4(\flow_control_config[31]_i_2_n_0 ),
        .I5(out[6]),
        .O(\flow_control_config[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \flow_control_config[31]_i_2 
       (.I0(out[3]),
        .I1(out[4]),
        .I2(out[7]),
        .I3(out[2]),
        .O(\flow_control_config[31]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[0] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[0]),
        .Q(\flow_control_config_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[10] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[10]),
        .Q(\flow_control_config_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[11] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[11]),
        .Q(\flow_control_config_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[12] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[12]),
        .Q(\flow_control_config_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[13] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[13]),
        .Q(\flow_control_config_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[14] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[14]),
        .Q(\flow_control_config_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[15] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[15]),
        .Q(\flow_control_config_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[16] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[16]),
        .Q(\flow_control_config_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[17] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[17]),
        .Q(\flow_control_config_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[18] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[18]),
        .Q(\flow_control_config_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[19] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[19]),
        .Q(\flow_control_config_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[1] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[1]),
        .Q(\flow_control_config_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[20] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[20]),
        .Q(\flow_control_config_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[21] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[21]),
        .Q(\flow_control_config_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[22] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[22]),
        .Q(\flow_control_config_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[23] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[23]),
        .Q(\flow_control_config_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[24] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[24]),
        .Q(\flow_control_config_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[25] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[25]),
        .Q(\flow_control_config_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[26] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[26]),
        .Q(\flow_control_config_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[27] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[27]),
        .Q(\flow_control_config_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[28] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[28]),
        .Q(\flow_control_config_reg_n_0_[28] ));
  FDPE #(
    .INIT(1'b1)) 
    \flow_control_config_reg[29] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .D(mgmt_wr_data[29]),
        .PRE(rst_i),
        .Q(\flow_control_config_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[2] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[2]),
        .Q(\flow_control_config_reg_n_0_[2] ));
  FDPE #(
    .INIT(1'b1)) 
    \flow_control_config_reg[30] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .D(mgmt_wr_data[30]),
        .PRE(rst_i),
        .Q(cfgTxRegData[0]));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[31] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[31]),
        .Q(\flow_control_config_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[3] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[3]),
        .Q(\flow_control_config_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[4] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[4]),
        .Q(\flow_control_config_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[5] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[5]),
        .Q(\flow_control_config_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[6] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[6]),
        .Q(\flow_control_config_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[7] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[7]),
        .Q(\flow_control_config_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[8] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[8]),
        .Q(\flow_control_config_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \flow_control_config_reg[9] 
       (.C(clk_i),
        .CE(\flow_control_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[9]),
        .Q(\flow_control_config_reg_n_0_[9] ));
  LUT1 #(
    .INIT(2'h1)) 
    \fragment_frame[0]_i_2 
       (.I0(fragment_frame_reg[0]),
        .O(\fragment_frame[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_15 ),
        .Q(fragment_frame_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[0]_i_1_n_0 ,\fragment_frame_reg[0]_i_1_n_1 ,\fragment_frame_reg[0]_i_1_n_2 ,\fragment_frame_reg[0]_i_1_n_3 ,\fragment_frame_reg[0]_i_1_n_4 ,\fragment_frame_reg[0]_i_1_n_5 ,\fragment_frame_reg[0]_i_1_n_6 ,\fragment_frame_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\fragment_frame_reg[0]_i_1_n_8 ,\fragment_frame_reg[0]_i_1_n_9 ,\fragment_frame_reg[0]_i_1_n_10 ,\fragment_frame_reg[0]_i_1_n_11 ,\fragment_frame_reg[0]_i_1_n_12 ,\fragment_frame_reg[0]_i_1_n_13 ,\fragment_frame_reg[0]_i_1_n_14 ,\fragment_frame_reg[0]_i_1_n_15 }),
        .S({fragment_frame_reg[7:1],\fragment_frame[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_13 ),
        .Q(fragment_frame_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_12 ),
        .Q(fragment_frame_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_11 ),
        .Q(fragment_frame_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_10 ),
        .Q(fragment_frame_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_9 ),
        .Q(fragment_frame_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_8 ),
        .Q(fragment_frame_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_15 ),
        .Q(fragment_frame_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[16]_i_1 
       (.CI(\fragment_frame_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[16]_i_1_n_0 ,\fragment_frame_reg[16]_i_1_n_1 ,\fragment_frame_reg[16]_i_1_n_2 ,\fragment_frame_reg[16]_i_1_n_3 ,\fragment_frame_reg[16]_i_1_n_4 ,\fragment_frame_reg[16]_i_1_n_5 ,\fragment_frame_reg[16]_i_1_n_6 ,\fragment_frame_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[16]_i_1_n_8 ,\fragment_frame_reg[16]_i_1_n_9 ,\fragment_frame_reg[16]_i_1_n_10 ,\fragment_frame_reg[16]_i_1_n_11 ,\fragment_frame_reg[16]_i_1_n_12 ,\fragment_frame_reg[16]_i_1_n_13 ,\fragment_frame_reg[16]_i_1_n_14 ,\fragment_frame_reg[16]_i_1_n_15 }),
        .S(fragment_frame_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_14 ),
        .Q(fragment_frame_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_13 ),
        .Q(fragment_frame_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_12 ),
        .Q(fragment_frame_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_14 ),
        .Q(fragment_frame_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_11 ),
        .Q(fragment_frame_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_10 ),
        .Q(fragment_frame_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_9 ),
        .Q(fragment_frame_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[16]_i_1_n_8 ),
        .Q(fragment_frame_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_15 ),
        .Q(fragment_frame_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[24]_i_1 
       (.CI(\fragment_frame_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[24]_i_1_n_0 ,\fragment_frame_reg[24]_i_1_n_1 ,\fragment_frame_reg[24]_i_1_n_2 ,\fragment_frame_reg[24]_i_1_n_3 ,\fragment_frame_reg[24]_i_1_n_4 ,\fragment_frame_reg[24]_i_1_n_5 ,\fragment_frame_reg[24]_i_1_n_6 ,\fragment_frame_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[24]_i_1_n_8 ,\fragment_frame_reg[24]_i_1_n_9 ,\fragment_frame_reg[24]_i_1_n_10 ,\fragment_frame_reg[24]_i_1_n_11 ,\fragment_frame_reg[24]_i_1_n_12 ,\fragment_frame_reg[24]_i_1_n_13 ,\fragment_frame_reg[24]_i_1_n_14 ,\fragment_frame_reg[24]_i_1_n_15 }),
        .S(fragment_frame_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_14 ),
        .Q(fragment_frame_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_13 ),
        .Q(fragment_frame_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_12 ),
        .Q(fragment_frame_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_11 ),
        .Q(fragment_frame_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_10 ),
        .Q(fragment_frame_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_13 ),
        .Q(fragment_frame_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_9 ),
        .Q(fragment_frame_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[24]_i_1_n_8 ),
        .Q(fragment_frame_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_15 ),
        .Q(fragment_frame_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[32]_i_1 
       (.CI(\fragment_frame_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[32]_i_1_n_0 ,\fragment_frame_reg[32]_i_1_n_1 ,\fragment_frame_reg[32]_i_1_n_2 ,\fragment_frame_reg[32]_i_1_n_3 ,\fragment_frame_reg[32]_i_1_n_4 ,\fragment_frame_reg[32]_i_1_n_5 ,\fragment_frame_reg[32]_i_1_n_6 ,\fragment_frame_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[32]_i_1_n_8 ,\fragment_frame_reg[32]_i_1_n_9 ,\fragment_frame_reg[32]_i_1_n_10 ,\fragment_frame_reg[32]_i_1_n_11 ,\fragment_frame_reg[32]_i_1_n_12 ,\fragment_frame_reg[32]_i_1_n_13 ,\fragment_frame_reg[32]_i_1_n_14 ,\fragment_frame_reg[32]_i_1_n_15 }),
        .S(fragment_frame_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_14 ),
        .Q(fragment_frame_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_13 ),
        .Q(fragment_frame_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_12 ),
        .Q(fragment_frame_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_11 ),
        .Q(fragment_frame_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_10 ),
        .Q(fragment_frame_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_9 ),
        .Q(fragment_frame_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[32]_i_1_n_8 ),
        .Q(fragment_frame_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_12 ),
        .Q(fragment_frame_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_15 ),
        .Q(fragment_frame_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[40]_i_1 
       (.CI(\fragment_frame_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[40]_i_1_n_0 ,\fragment_frame_reg[40]_i_1_n_1 ,\fragment_frame_reg[40]_i_1_n_2 ,\fragment_frame_reg[40]_i_1_n_3 ,\fragment_frame_reg[40]_i_1_n_4 ,\fragment_frame_reg[40]_i_1_n_5 ,\fragment_frame_reg[40]_i_1_n_6 ,\fragment_frame_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[40]_i_1_n_8 ,\fragment_frame_reg[40]_i_1_n_9 ,\fragment_frame_reg[40]_i_1_n_10 ,\fragment_frame_reg[40]_i_1_n_11 ,\fragment_frame_reg[40]_i_1_n_12 ,\fragment_frame_reg[40]_i_1_n_13 ,\fragment_frame_reg[40]_i_1_n_14 ,\fragment_frame_reg[40]_i_1_n_15 }),
        .S(fragment_frame_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_14 ),
        .Q(fragment_frame_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_13 ),
        .Q(fragment_frame_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_12 ),
        .Q(fragment_frame_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_11 ),
        .Q(fragment_frame_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_10 ),
        .Q(fragment_frame_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_9 ),
        .Q(fragment_frame_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[40]_i_1_n_8 ),
        .Q(fragment_frame_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_15 ),
        .Q(fragment_frame_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[48]_i_1 
       (.CI(\fragment_frame_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[48]_i_1_n_0 ,\fragment_frame_reg[48]_i_1_n_1 ,\fragment_frame_reg[48]_i_1_n_2 ,\fragment_frame_reg[48]_i_1_n_3 ,\fragment_frame_reg[48]_i_1_n_4 ,\fragment_frame_reg[48]_i_1_n_5 ,\fragment_frame_reg[48]_i_1_n_6 ,\fragment_frame_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[48]_i_1_n_8 ,\fragment_frame_reg[48]_i_1_n_9 ,\fragment_frame_reg[48]_i_1_n_10 ,\fragment_frame_reg[48]_i_1_n_11 ,\fragment_frame_reg[48]_i_1_n_12 ,\fragment_frame_reg[48]_i_1_n_13 ,\fragment_frame_reg[48]_i_1_n_14 ,\fragment_frame_reg[48]_i_1_n_15 }),
        .S(fragment_frame_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_14 ),
        .Q(fragment_frame_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_11 ),
        .Q(fragment_frame_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_13 ),
        .Q(fragment_frame_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_12 ),
        .Q(fragment_frame_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_11 ),
        .Q(fragment_frame_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_10 ),
        .Q(fragment_frame_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_9 ),
        .Q(fragment_frame_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[48]_i_1_n_8 ),
        .Q(fragment_frame_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_15 ),
        .Q(fragment_frame_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[56]_i_1 
       (.CI(\fragment_frame_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_fragment_frame_reg[56]_i_1_CO_UNCONNECTED [7],\fragment_frame_reg[56]_i_1_n_1 ,\fragment_frame_reg[56]_i_1_n_2 ,\fragment_frame_reg[56]_i_1_n_3 ,\fragment_frame_reg[56]_i_1_n_4 ,\fragment_frame_reg[56]_i_1_n_5 ,\fragment_frame_reg[56]_i_1_n_6 ,\fragment_frame_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[56]_i_1_n_8 ,\fragment_frame_reg[56]_i_1_n_9 ,\fragment_frame_reg[56]_i_1_n_10 ,\fragment_frame_reg[56]_i_1_n_11 ,\fragment_frame_reg[56]_i_1_n_12 ,\fragment_frame_reg[56]_i_1_n_13 ,\fragment_frame_reg[56]_i_1_n_14 ,\fragment_frame_reg[56]_i_1_n_15 }),
        .S(fragment_frame_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_14 ),
        .Q(fragment_frame_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_13 ),
        .Q(fragment_frame_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_12 ),
        .Q(fragment_frame_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_10 ),
        .Q(fragment_frame_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_11 ),
        .Q(fragment_frame_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_10 ),
        .Q(fragment_frame_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_9 ),
        .Q(fragment_frame_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[56]_i_1_n_8 ),
        .Q(fragment_frame_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_9 ),
        .Q(fragment_frame_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[0]_i_1_n_8 ),
        .Q(fragment_frame_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_15 ),
        .Q(fragment_frame_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \fragment_frame_reg[8]_i_1 
       (.CI(\fragment_frame_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\fragment_frame_reg[8]_i_1_n_0 ,\fragment_frame_reg[8]_i_1_n_1 ,\fragment_frame_reg[8]_i_1_n_2 ,\fragment_frame_reg[8]_i_1_n_3 ,\fragment_frame_reg[8]_i_1_n_4 ,\fragment_frame_reg[8]_i_1_n_5 ,\fragment_frame_reg[8]_i_1_n_6 ,\fragment_frame_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\fragment_frame_reg[8]_i_1_n_8 ,\fragment_frame_reg[8]_i_1_n_9 ,\fragment_frame_reg[8]_i_1_n_10 ,\fragment_frame_reg[8]_i_1_n_11 ,\fragment_frame_reg[8]_i_1_n_12 ,\fragment_frame_reg[8]_i_1_n_13 ,\fragment_frame_reg[8]_i_1_n_14 ,\fragment_frame_reg[8]_i_1_n_15 }),
        .S(fragment_frame_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \fragment_frame_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[17]),
        .CLR(rst_i),
        .D(\fragment_frame_reg[8]_i_1_n_14 ),
        .Q(fragment_frame_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_1024_max_good[0]_i_2 
       (.I0(frame_1024_max_good_reg[0]),
        .O(\frame_1024_max_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[0]_i_1_n_0 ,\frame_1024_max_good_reg[0]_i_1_n_1 ,\frame_1024_max_good_reg[0]_i_1_n_2 ,\frame_1024_max_good_reg[0]_i_1_n_3 ,\frame_1024_max_good_reg[0]_i_1_n_4 ,\frame_1024_max_good_reg[0]_i_1_n_5 ,\frame_1024_max_good_reg[0]_i_1_n_6 ,\frame_1024_max_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_1024_max_good_reg[0]_i_1_n_8 ,\frame_1024_max_good_reg[0]_i_1_n_9 ,\frame_1024_max_good_reg[0]_i_1_n_10 ,\frame_1024_max_good_reg[0]_i_1_n_11 ,\frame_1024_max_good_reg[0]_i_1_n_12 ,\frame_1024_max_good_reg[0]_i_1_n_13 ,\frame_1024_max_good_reg[0]_i_1_n_14 ,\frame_1024_max_good_reg[0]_i_1_n_15 }),
        .S({frame_1024_max_good_reg[7:1],\frame_1024_max_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[16]_i_1 
       (.CI(\frame_1024_max_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[16]_i_1_n_0 ,\frame_1024_max_good_reg[16]_i_1_n_1 ,\frame_1024_max_good_reg[16]_i_1_n_2 ,\frame_1024_max_good_reg[16]_i_1_n_3 ,\frame_1024_max_good_reg[16]_i_1_n_4 ,\frame_1024_max_good_reg[16]_i_1_n_5 ,\frame_1024_max_good_reg[16]_i_1_n_6 ,\frame_1024_max_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[16]_i_1_n_8 ,\frame_1024_max_good_reg[16]_i_1_n_9 ,\frame_1024_max_good_reg[16]_i_1_n_10 ,\frame_1024_max_good_reg[16]_i_1_n_11 ,\frame_1024_max_good_reg[16]_i_1_n_12 ,\frame_1024_max_good_reg[16]_i_1_n_13 ,\frame_1024_max_good_reg[16]_i_1_n_14 ,\frame_1024_max_good_reg[16]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[16]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[24]_i_1 
       (.CI(\frame_1024_max_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[24]_i_1_n_0 ,\frame_1024_max_good_reg[24]_i_1_n_1 ,\frame_1024_max_good_reg[24]_i_1_n_2 ,\frame_1024_max_good_reg[24]_i_1_n_3 ,\frame_1024_max_good_reg[24]_i_1_n_4 ,\frame_1024_max_good_reg[24]_i_1_n_5 ,\frame_1024_max_good_reg[24]_i_1_n_6 ,\frame_1024_max_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[24]_i_1_n_8 ,\frame_1024_max_good_reg[24]_i_1_n_9 ,\frame_1024_max_good_reg[24]_i_1_n_10 ,\frame_1024_max_good_reg[24]_i_1_n_11 ,\frame_1024_max_good_reg[24]_i_1_n_12 ,\frame_1024_max_good_reg[24]_i_1_n_13 ,\frame_1024_max_good_reg[24]_i_1_n_14 ,\frame_1024_max_good_reg[24]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[24]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[32]_i_1 
       (.CI(\frame_1024_max_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[32]_i_1_n_0 ,\frame_1024_max_good_reg[32]_i_1_n_1 ,\frame_1024_max_good_reg[32]_i_1_n_2 ,\frame_1024_max_good_reg[32]_i_1_n_3 ,\frame_1024_max_good_reg[32]_i_1_n_4 ,\frame_1024_max_good_reg[32]_i_1_n_5 ,\frame_1024_max_good_reg[32]_i_1_n_6 ,\frame_1024_max_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[32]_i_1_n_8 ,\frame_1024_max_good_reg[32]_i_1_n_9 ,\frame_1024_max_good_reg[32]_i_1_n_10 ,\frame_1024_max_good_reg[32]_i_1_n_11 ,\frame_1024_max_good_reg[32]_i_1_n_12 ,\frame_1024_max_good_reg[32]_i_1_n_13 ,\frame_1024_max_good_reg[32]_i_1_n_14 ,\frame_1024_max_good_reg[32]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[32]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[40]_i_1 
       (.CI(\frame_1024_max_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[40]_i_1_n_0 ,\frame_1024_max_good_reg[40]_i_1_n_1 ,\frame_1024_max_good_reg[40]_i_1_n_2 ,\frame_1024_max_good_reg[40]_i_1_n_3 ,\frame_1024_max_good_reg[40]_i_1_n_4 ,\frame_1024_max_good_reg[40]_i_1_n_5 ,\frame_1024_max_good_reg[40]_i_1_n_6 ,\frame_1024_max_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[40]_i_1_n_8 ,\frame_1024_max_good_reg[40]_i_1_n_9 ,\frame_1024_max_good_reg[40]_i_1_n_10 ,\frame_1024_max_good_reg[40]_i_1_n_11 ,\frame_1024_max_good_reg[40]_i_1_n_12 ,\frame_1024_max_good_reg[40]_i_1_n_13 ,\frame_1024_max_good_reg[40]_i_1_n_14 ,\frame_1024_max_good_reg[40]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[40]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[48]_i_1 
       (.CI(\frame_1024_max_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[48]_i_1_n_0 ,\frame_1024_max_good_reg[48]_i_1_n_1 ,\frame_1024_max_good_reg[48]_i_1_n_2 ,\frame_1024_max_good_reg[48]_i_1_n_3 ,\frame_1024_max_good_reg[48]_i_1_n_4 ,\frame_1024_max_good_reg[48]_i_1_n_5 ,\frame_1024_max_good_reg[48]_i_1_n_6 ,\frame_1024_max_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[48]_i_1_n_8 ,\frame_1024_max_good_reg[48]_i_1_n_9 ,\frame_1024_max_good_reg[48]_i_1_n_10 ,\frame_1024_max_good_reg[48]_i_1_n_11 ,\frame_1024_max_good_reg[48]_i_1_n_12 ,\frame_1024_max_good_reg[48]_i_1_n_13 ,\frame_1024_max_good_reg[48]_i_1_n_14 ,\frame_1024_max_good_reg[48]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[48]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[56]_i_1 
       (.CI(\frame_1024_max_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_1024_max_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_1024_max_good_reg[56]_i_1_n_1 ,\frame_1024_max_good_reg[56]_i_1_n_2 ,\frame_1024_max_good_reg[56]_i_1_n_3 ,\frame_1024_max_good_reg[56]_i_1_n_4 ,\frame_1024_max_good_reg[56]_i_1_n_5 ,\frame_1024_max_good_reg[56]_i_1_n_6 ,\frame_1024_max_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[56]_i_1_n_8 ,\frame_1024_max_good_reg[56]_i_1_n_9 ,\frame_1024_max_good_reg[56]_i_1_n_10 ,\frame_1024_max_good_reg[56]_i_1_n_11 ,\frame_1024_max_good_reg[56]_i_1_n_12 ,\frame_1024_max_good_reg[56]_i_1_n_13 ,\frame_1024_max_good_reg[56]_i_1_n_14 ,\frame_1024_max_good_reg[56]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_13 ),
        .Q(frame_1024_max_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_12 ),
        .Q(frame_1024_max_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_11 ),
        .Q(frame_1024_max_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_10 ),
        .Q(frame_1024_max_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[56]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_9 ),
        .Q(frame_1024_max_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[0]_i_1_n_8 ),
        .Q(frame_1024_max_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_15 ),
        .Q(frame_1024_max_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_good_reg[8]_i_1 
       (.CI(\frame_1024_max_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_good_reg[8]_i_1_n_0 ,\frame_1024_max_good_reg[8]_i_1_n_1 ,\frame_1024_max_good_reg[8]_i_1_n_2 ,\frame_1024_max_good_reg[8]_i_1_n_3 ,\frame_1024_max_good_reg[8]_i_1_n_4 ,\frame_1024_max_good_reg[8]_i_1_n_5 ,\frame_1024_max_good_reg[8]_i_1_n_6 ,\frame_1024_max_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_good_reg[8]_i_1_n_8 ,\frame_1024_max_good_reg[8]_i_1_n_9 ,\frame_1024_max_good_reg[8]_i_1_n_10 ,\frame_1024_max_good_reg[8]_i_1_n_11 ,\frame_1024_max_good_reg[8]_i_1_n_12 ,\frame_1024_max_good_reg[8]_i_1_n_13 ,\frame_1024_max_good_reg[8]_i_1_n_14 ,\frame_1024_max_good_reg[8]_i_1_n_15 }),
        .S(frame_1024_max_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_1024_max_good_reg[8]_i_1_n_14 ),
        .Q(frame_1024_max_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_1024_max_transed[0]_i_2 
       (.I0(frame_1024_max_transed_reg[0]),
        .O(\frame_1024_max_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[0]_i_1_n_0 ,\frame_1024_max_transed_reg[0]_i_1_n_1 ,\frame_1024_max_transed_reg[0]_i_1_n_2 ,\frame_1024_max_transed_reg[0]_i_1_n_3 ,\frame_1024_max_transed_reg[0]_i_1_n_4 ,\frame_1024_max_transed_reg[0]_i_1_n_5 ,\frame_1024_max_transed_reg[0]_i_1_n_6 ,\frame_1024_max_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_1024_max_transed_reg[0]_i_1_n_8 ,\frame_1024_max_transed_reg[0]_i_1_n_9 ,\frame_1024_max_transed_reg[0]_i_1_n_10 ,\frame_1024_max_transed_reg[0]_i_1_n_11 ,\frame_1024_max_transed_reg[0]_i_1_n_12 ,\frame_1024_max_transed_reg[0]_i_1_n_13 ,\frame_1024_max_transed_reg[0]_i_1_n_14 ,\frame_1024_max_transed_reg[0]_i_1_n_15 }),
        .S({frame_1024_max_transed_reg[7:1],\frame_1024_max_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[16]_i_1 
       (.CI(\frame_1024_max_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[16]_i_1_n_0 ,\frame_1024_max_transed_reg[16]_i_1_n_1 ,\frame_1024_max_transed_reg[16]_i_1_n_2 ,\frame_1024_max_transed_reg[16]_i_1_n_3 ,\frame_1024_max_transed_reg[16]_i_1_n_4 ,\frame_1024_max_transed_reg[16]_i_1_n_5 ,\frame_1024_max_transed_reg[16]_i_1_n_6 ,\frame_1024_max_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[16]_i_1_n_8 ,\frame_1024_max_transed_reg[16]_i_1_n_9 ,\frame_1024_max_transed_reg[16]_i_1_n_10 ,\frame_1024_max_transed_reg[16]_i_1_n_11 ,\frame_1024_max_transed_reg[16]_i_1_n_12 ,\frame_1024_max_transed_reg[16]_i_1_n_13 ,\frame_1024_max_transed_reg[16]_i_1_n_14 ,\frame_1024_max_transed_reg[16]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[16]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[24]_i_1 
       (.CI(\frame_1024_max_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[24]_i_1_n_0 ,\frame_1024_max_transed_reg[24]_i_1_n_1 ,\frame_1024_max_transed_reg[24]_i_1_n_2 ,\frame_1024_max_transed_reg[24]_i_1_n_3 ,\frame_1024_max_transed_reg[24]_i_1_n_4 ,\frame_1024_max_transed_reg[24]_i_1_n_5 ,\frame_1024_max_transed_reg[24]_i_1_n_6 ,\frame_1024_max_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[24]_i_1_n_8 ,\frame_1024_max_transed_reg[24]_i_1_n_9 ,\frame_1024_max_transed_reg[24]_i_1_n_10 ,\frame_1024_max_transed_reg[24]_i_1_n_11 ,\frame_1024_max_transed_reg[24]_i_1_n_12 ,\frame_1024_max_transed_reg[24]_i_1_n_13 ,\frame_1024_max_transed_reg[24]_i_1_n_14 ,\frame_1024_max_transed_reg[24]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[24]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[32]_i_1 
       (.CI(\frame_1024_max_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[32]_i_1_n_0 ,\frame_1024_max_transed_reg[32]_i_1_n_1 ,\frame_1024_max_transed_reg[32]_i_1_n_2 ,\frame_1024_max_transed_reg[32]_i_1_n_3 ,\frame_1024_max_transed_reg[32]_i_1_n_4 ,\frame_1024_max_transed_reg[32]_i_1_n_5 ,\frame_1024_max_transed_reg[32]_i_1_n_6 ,\frame_1024_max_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[32]_i_1_n_8 ,\frame_1024_max_transed_reg[32]_i_1_n_9 ,\frame_1024_max_transed_reg[32]_i_1_n_10 ,\frame_1024_max_transed_reg[32]_i_1_n_11 ,\frame_1024_max_transed_reg[32]_i_1_n_12 ,\frame_1024_max_transed_reg[32]_i_1_n_13 ,\frame_1024_max_transed_reg[32]_i_1_n_14 ,\frame_1024_max_transed_reg[32]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[32]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[40]_i_1 
       (.CI(\frame_1024_max_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[40]_i_1_n_0 ,\frame_1024_max_transed_reg[40]_i_1_n_1 ,\frame_1024_max_transed_reg[40]_i_1_n_2 ,\frame_1024_max_transed_reg[40]_i_1_n_3 ,\frame_1024_max_transed_reg[40]_i_1_n_4 ,\frame_1024_max_transed_reg[40]_i_1_n_5 ,\frame_1024_max_transed_reg[40]_i_1_n_6 ,\frame_1024_max_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[40]_i_1_n_8 ,\frame_1024_max_transed_reg[40]_i_1_n_9 ,\frame_1024_max_transed_reg[40]_i_1_n_10 ,\frame_1024_max_transed_reg[40]_i_1_n_11 ,\frame_1024_max_transed_reg[40]_i_1_n_12 ,\frame_1024_max_transed_reg[40]_i_1_n_13 ,\frame_1024_max_transed_reg[40]_i_1_n_14 ,\frame_1024_max_transed_reg[40]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[40]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[48]_i_1 
       (.CI(\frame_1024_max_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[48]_i_1_n_0 ,\frame_1024_max_transed_reg[48]_i_1_n_1 ,\frame_1024_max_transed_reg[48]_i_1_n_2 ,\frame_1024_max_transed_reg[48]_i_1_n_3 ,\frame_1024_max_transed_reg[48]_i_1_n_4 ,\frame_1024_max_transed_reg[48]_i_1_n_5 ,\frame_1024_max_transed_reg[48]_i_1_n_6 ,\frame_1024_max_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[48]_i_1_n_8 ,\frame_1024_max_transed_reg[48]_i_1_n_9 ,\frame_1024_max_transed_reg[48]_i_1_n_10 ,\frame_1024_max_transed_reg[48]_i_1_n_11 ,\frame_1024_max_transed_reg[48]_i_1_n_12 ,\frame_1024_max_transed_reg[48]_i_1_n_13 ,\frame_1024_max_transed_reg[48]_i_1_n_14 ,\frame_1024_max_transed_reg[48]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[48]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[56]_i_1 
       (.CI(\frame_1024_max_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_1024_max_transed_reg[56]_i_1_CO_UNCONNECTED [7],\frame_1024_max_transed_reg[56]_i_1_n_1 ,\frame_1024_max_transed_reg[56]_i_1_n_2 ,\frame_1024_max_transed_reg[56]_i_1_n_3 ,\frame_1024_max_transed_reg[56]_i_1_n_4 ,\frame_1024_max_transed_reg[56]_i_1_n_5 ,\frame_1024_max_transed_reg[56]_i_1_n_6 ,\frame_1024_max_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[56]_i_1_n_8 ,\frame_1024_max_transed_reg[56]_i_1_n_9 ,\frame_1024_max_transed_reg[56]_i_1_n_10 ,\frame_1024_max_transed_reg[56]_i_1_n_11 ,\frame_1024_max_transed_reg[56]_i_1_n_12 ,\frame_1024_max_transed_reg[56]_i_1_n_13 ,\frame_1024_max_transed_reg[56]_i_1_n_14 ,\frame_1024_max_transed_reg[56]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_13 ),
        .Q(frame_1024_max_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_12 ),
        .Q(frame_1024_max_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_11 ),
        .Q(frame_1024_max_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_10 ),
        .Q(frame_1024_max_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[56]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_9 ),
        .Q(frame_1024_max_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[0]_i_1_n_8 ),
        .Q(frame_1024_max_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_15 ),
        .Q(frame_1024_max_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_1024_max_transed_reg[8]_i_1 
       (.CI(\frame_1024_max_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_1024_max_transed_reg[8]_i_1_n_0 ,\frame_1024_max_transed_reg[8]_i_1_n_1 ,\frame_1024_max_transed_reg[8]_i_1_n_2 ,\frame_1024_max_transed_reg[8]_i_1_n_3 ,\frame_1024_max_transed_reg[8]_i_1_n_4 ,\frame_1024_max_transed_reg[8]_i_1_n_5 ,\frame_1024_max_transed_reg[8]_i_1_n_6 ,\frame_1024_max_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_1024_max_transed_reg[8]_i_1_n_8 ,\frame_1024_max_transed_reg[8]_i_1_n_9 ,\frame_1024_max_transed_reg[8]_i_1_n_10 ,\frame_1024_max_transed_reg[8]_i_1_n_11 ,\frame_1024_max_transed_reg[8]_i_1_n_12 ,\frame_1024_max_transed_reg[8]_i_1_n_13 ,\frame_1024_max_transed_reg[8]_i_1_n_14 ,\frame_1024_max_transed_reg[8]_i_1_n_15 }),
        .S(frame_1024_max_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_1024_max_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[11]),
        .CLR(rst_i),
        .D(\frame_1024_max_transed_reg[8]_i_1_n_14 ),
        .Q(frame_1024_max_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_128_255_good[0]_i_2 
       (.I0(frame_128_255_good_reg[0]),
        .O(\frame_128_255_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[0]_i_1_n_0 ,\frame_128_255_good_reg[0]_i_1_n_1 ,\frame_128_255_good_reg[0]_i_1_n_2 ,\frame_128_255_good_reg[0]_i_1_n_3 ,\frame_128_255_good_reg[0]_i_1_n_4 ,\frame_128_255_good_reg[0]_i_1_n_5 ,\frame_128_255_good_reg[0]_i_1_n_6 ,\frame_128_255_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_128_255_good_reg[0]_i_1_n_8 ,\frame_128_255_good_reg[0]_i_1_n_9 ,\frame_128_255_good_reg[0]_i_1_n_10 ,\frame_128_255_good_reg[0]_i_1_n_11 ,\frame_128_255_good_reg[0]_i_1_n_12 ,\frame_128_255_good_reg[0]_i_1_n_13 ,\frame_128_255_good_reg[0]_i_1_n_14 ,\frame_128_255_good_reg[0]_i_1_n_15 }),
        .S({frame_128_255_good_reg[7:1],\frame_128_255_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[16]_i_1 
       (.CI(\frame_128_255_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[16]_i_1_n_0 ,\frame_128_255_good_reg[16]_i_1_n_1 ,\frame_128_255_good_reg[16]_i_1_n_2 ,\frame_128_255_good_reg[16]_i_1_n_3 ,\frame_128_255_good_reg[16]_i_1_n_4 ,\frame_128_255_good_reg[16]_i_1_n_5 ,\frame_128_255_good_reg[16]_i_1_n_6 ,\frame_128_255_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[16]_i_1_n_8 ,\frame_128_255_good_reg[16]_i_1_n_9 ,\frame_128_255_good_reg[16]_i_1_n_10 ,\frame_128_255_good_reg[16]_i_1_n_11 ,\frame_128_255_good_reg[16]_i_1_n_12 ,\frame_128_255_good_reg[16]_i_1_n_13 ,\frame_128_255_good_reg[16]_i_1_n_14 ,\frame_128_255_good_reg[16]_i_1_n_15 }),
        .S(frame_128_255_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[16]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[24]_i_1 
       (.CI(\frame_128_255_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[24]_i_1_n_0 ,\frame_128_255_good_reg[24]_i_1_n_1 ,\frame_128_255_good_reg[24]_i_1_n_2 ,\frame_128_255_good_reg[24]_i_1_n_3 ,\frame_128_255_good_reg[24]_i_1_n_4 ,\frame_128_255_good_reg[24]_i_1_n_5 ,\frame_128_255_good_reg[24]_i_1_n_6 ,\frame_128_255_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[24]_i_1_n_8 ,\frame_128_255_good_reg[24]_i_1_n_9 ,\frame_128_255_good_reg[24]_i_1_n_10 ,\frame_128_255_good_reg[24]_i_1_n_11 ,\frame_128_255_good_reg[24]_i_1_n_12 ,\frame_128_255_good_reg[24]_i_1_n_13 ,\frame_128_255_good_reg[24]_i_1_n_14 ,\frame_128_255_good_reg[24]_i_1_n_15 }),
        .S(frame_128_255_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[24]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[32]_i_1 
       (.CI(\frame_128_255_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[32]_i_1_n_0 ,\frame_128_255_good_reg[32]_i_1_n_1 ,\frame_128_255_good_reg[32]_i_1_n_2 ,\frame_128_255_good_reg[32]_i_1_n_3 ,\frame_128_255_good_reg[32]_i_1_n_4 ,\frame_128_255_good_reg[32]_i_1_n_5 ,\frame_128_255_good_reg[32]_i_1_n_6 ,\frame_128_255_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[32]_i_1_n_8 ,\frame_128_255_good_reg[32]_i_1_n_9 ,\frame_128_255_good_reg[32]_i_1_n_10 ,\frame_128_255_good_reg[32]_i_1_n_11 ,\frame_128_255_good_reg[32]_i_1_n_12 ,\frame_128_255_good_reg[32]_i_1_n_13 ,\frame_128_255_good_reg[32]_i_1_n_14 ,\frame_128_255_good_reg[32]_i_1_n_15 }),
        .S(frame_128_255_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[32]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[40]_i_1 
       (.CI(\frame_128_255_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[40]_i_1_n_0 ,\frame_128_255_good_reg[40]_i_1_n_1 ,\frame_128_255_good_reg[40]_i_1_n_2 ,\frame_128_255_good_reg[40]_i_1_n_3 ,\frame_128_255_good_reg[40]_i_1_n_4 ,\frame_128_255_good_reg[40]_i_1_n_5 ,\frame_128_255_good_reg[40]_i_1_n_6 ,\frame_128_255_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[40]_i_1_n_8 ,\frame_128_255_good_reg[40]_i_1_n_9 ,\frame_128_255_good_reg[40]_i_1_n_10 ,\frame_128_255_good_reg[40]_i_1_n_11 ,\frame_128_255_good_reg[40]_i_1_n_12 ,\frame_128_255_good_reg[40]_i_1_n_13 ,\frame_128_255_good_reg[40]_i_1_n_14 ,\frame_128_255_good_reg[40]_i_1_n_15 }),
        .S(frame_128_255_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[40]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[48]_i_1 
       (.CI(\frame_128_255_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[48]_i_1_n_0 ,\frame_128_255_good_reg[48]_i_1_n_1 ,\frame_128_255_good_reg[48]_i_1_n_2 ,\frame_128_255_good_reg[48]_i_1_n_3 ,\frame_128_255_good_reg[48]_i_1_n_4 ,\frame_128_255_good_reg[48]_i_1_n_5 ,\frame_128_255_good_reg[48]_i_1_n_6 ,\frame_128_255_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[48]_i_1_n_8 ,\frame_128_255_good_reg[48]_i_1_n_9 ,\frame_128_255_good_reg[48]_i_1_n_10 ,\frame_128_255_good_reg[48]_i_1_n_11 ,\frame_128_255_good_reg[48]_i_1_n_12 ,\frame_128_255_good_reg[48]_i_1_n_13 ,\frame_128_255_good_reg[48]_i_1_n_14 ,\frame_128_255_good_reg[48]_i_1_n_15 }),
        .S(frame_128_255_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[48]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[56]_i_1 
       (.CI(\frame_128_255_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_128_255_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_128_255_good_reg[56]_i_1_n_1 ,\frame_128_255_good_reg[56]_i_1_n_2 ,\frame_128_255_good_reg[56]_i_1_n_3 ,\frame_128_255_good_reg[56]_i_1_n_4 ,\frame_128_255_good_reg[56]_i_1_n_5 ,\frame_128_255_good_reg[56]_i_1_n_6 ,\frame_128_255_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[56]_i_1_n_8 ,\frame_128_255_good_reg[56]_i_1_n_9 ,\frame_128_255_good_reg[56]_i_1_n_10 ,\frame_128_255_good_reg[56]_i_1_n_11 ,\frame_128_255_good_reg[56]_i_1_n_12 ,\frame_128_255_good_reg[56]_i_1_n_13 ,\frame_128_255_good_reg[56]_i_1_n_14 ,\frame_128_255_good_reg[56]_i_1_n_15 }),
        .S(frame_128_255_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_13 ),
        .Q(frame_128_255_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_12 ),
        .Q(frame_128_255_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_11 ),
        .Q(frame_128_255_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_10 ),
        .Q(frame_128_255_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[56]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_9 ),
        .Q(frame_128_255_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[0]_i_1_n_8 ),
        .Q(frame_128_255_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_15 ),
        .Q(frame_128_255_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_good_reg[8]_i_1 
       (.CI(\frame_128_255_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_good_reg[8]_i_1_n_0 ,\frame_128_255_good_reg[8]_i_1_n_1 ,\frame_128_255_good_reg[8]_i_1_n_2 ,\frame_128_255_good_reg[8]_i_1_n_3 ,\frame_128_255_good_reg[8]_i_1_n_4 ,\frame_128_255_good_reg[8]_i_1_n_5 ,\frame_128_255_good_reg[8]_i_1_n_6 ,\frame_128_255_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_good_reg[8]_i_1_n_8 ,\frame_128_255_good_reg[8]_i_1_n_9 ,\frame_128_255_good_reg[8]_i_1_n_10 ,\frame_128_255_good_reg[8]_i_1_n_11 ,\frame_128_255_good_reg[8]_i_1_n_12 ,\frame_128_255_good_reg[8]_i_1_n_13 ,\frame_128_255_good_reg[8]_i_1_n_14 ,\frame_128_255_good_reg[8]_i_1_n_15 }),
        .S(frame_128_255_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_128_255_good_reg[8]_i_1_n_14 ),
        .Q(frame_128_255_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_128_255_transed[0]_i_2 
       (.I0(frame_128_255_transed_reg[0]),
        .O(\frame_128_255_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[0]_i_1_n_0 ,\frame_128_255_transed_reg[0]_i_1_n_1 ,\frame_128_255_transed_reg[0]_i_1_n_2 ,\frame_128_255_transed_reg[0]_i_1_n_3 ,\frame_128_255_transed_reg[0]_i_1_n_4 ,\frame_128_255_transed_reg[0]_i_1_n_5 ,\frame_128_255_transed_reg[0]_i_1_n_6 ,\frame_128_255_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_128_255_transed_reg[0]_i_1_n_8 ,\frame_128_255_transed_reg[0]_i_1_n_9 ,\frame_128_255_transed_reg[0]_i_1_n_10 ,\frame_128_255_transed_reg[0]_i_1_n_11 ,\frame_128_255_transed_reg[0]_i_1_n_12 ,\frame_128_255_transed_reg[0]_i_1_n_13 ,\frame_128_255_transed_reg[0]_i_1_n_14 ,\frame_128_255_transed_reg[0]_i_1_n_15 }),
        .S({frame_128_255_transed_reg[7:1],\frame_128_255_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[16]_i_1 
       (.CI(\frame_128_255_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[16]_i_1_n_0 ,\frame_128_255_transed_reg[16]_i_1_n_1 ,\frame_128_255_transed_reg[16]_i_1_n_2 ,\frame_128_255_transed_reg[16]_i_1_n_3 ,\frame_128_255_transed_reg[16]_i_1_n_4 ,\frame_128_255_transed_reg[16]_i_1_n_5 ,\frame_128_255_transed_reg[16]_i_1_n_6 ,\frame_128_255_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[16]_i_1_n_8 ,\frame_128_255_transed_reg[16]_i_1_n_9 ,\frame_128_255_transed_reg[16]_i_1_n_10 ,\frame_128_255_transed_reg[16]_i_1_n_11 ,\frame_128_255_transed_reg[16]_i_1_n_12 ,\frame_128_255_transed_reg[16]_i_1_n_13 ,\frame_128_255_transed_reg[16]_i_1_n_14 ,\frame_128_255_transed_reg[16]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[16]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[24]_i_1 
       (.CI(\frame_128_255_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[24]_i_1_n_0 ,\frame_128_255_transed_reg[24]_i_1_n_1 ,\frame_128_255_transed_reg[24]_i_1_n_2 ,\frame_128_255_transed_reg[24]_i_1_n_3 ,\frame_128_255_transed_reg[24]_i_1_n_4 ,\frame_128_255_transed_reg[24]_i_1_n_5 ,\frame_128_255_transed_reg[24]_i_1_n_6 ,\frame_128_255_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[24]_i_1_n_8 ,\frame_128_255_transed_reg[24]_i_1_n_9 ,\frame_128_255_transed_reg[24]_i_1_n_10 ,\frame_128_255_transed_reg[24]_i_1_n_11 ,\frame_128_255_transed_reg[24]_i_1_n_12 ,\frame_128_255_transed_reg[24]_i_1_n_13 ,\frame_128_255_transed_reg[24]_i_1_n_14 ,\frame_128_255_transed_reg[24]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[24]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[32]_i_1 
       (.CI(\frame_128_255_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[32]_i_1_n_0 ,\frame_128_255_transed_reg[32]_i_1_n_1 ,\frame_128_255_transed_reg[32]_i_1_n_2 ,\frame_128_255_transed_reg[32]_i_1_n_3 ,\frame_128_255_transed_reg[32]_i_1_n_4 ,\frame_128_255_transed_reg[32]_i_1_n_5 ,\frame_128_255_transed_reg[32]_i_1_n_6 ,\frame_128_255_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[32]_i_1_n_8 ,\frame_128_255_transed_reg[32]_i_1_n_9 ,\frame_128_255_transed_reg[32]_i_1_n_10 ,\frame_128_255_transed_reg[32]_i_1_n_11 ,\frame_128_255_transed_reg[32]_i_1_n_12 ,\frame_128_255_transed_reg[32]_i_1_n_13 ,\frame_128_255_transed_reg[32]_i_1_n_14 ,\frame_128_255_transed_reg[32]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[32]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[40]_i_1 
       (.CI(\frame_128_255_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[40]_i_1_n_0 ,\frame_128_255_transed_reg[40]_i_1_n_1 ,\frame_128_255_transed_reg[40]_i_1_n_2 ,\frame_128_255_transed_reg[40]_i_1_n_3 ,\frame_128_255_transed_reg[40]_i_1_n_4 ,\frame_128_255_transed_reg[40]_i_1_n_5 ,\frame_128_255_transed_reg[40]_i_1_n_6 ,\frame_128_255_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[40]_i_1_n_8 ,\frame_128_255_transed_reg[40]_i_1_n_9 ,\frame_128_255_transed_reg[40]_i_1_n_10 ,\frame_128_255_transed_reg[40]_i_1_n_11 ,\frame_128_255_transed_reg[40]_i_1_n_12 ,\frame_128_255_transed_reg[40]_i_1_n_13 ,\frame_128_255_transed_reg[40]_i_1_n_14 ,\frame_128_255_transed_reg[40]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[40]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[48]_i_1 
       (.CI(\frame_128_255_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[48]_i_1_n_0 ,\frame_128_255_transed_reg[48]_i_1_n_1 ,\frame_128_255_transed_reg[48]_i_1_n_2 ,\frame_128_255_transed_reg[48]_i_1_n_3 ,\frame_128_255_transed_reg[48]_i_1_n_4 ,\frame_128_255_transed_reg[48]_i_1_n_5 ,\frame_128_255_transed_reg[48]_i_1_n_6 ,\frame_128_255_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[48]_i_1_n_8 ,\frame_128_255_transed_reg[48]_i_1_n_9 ,\frame_128_255_transed_reg[48]_i_1_n_10 ,\frame_128_255_transed_reg[48]_i_1_n_11 ,\frame_128_255_transed_reg[48]_i_1_n_12 ,\frame_128_255_transed_reg[48]_i_1_n_13 ,\frame_128_255_transed_reg[48]_i_1_n_14 ,\frame_128_255_transed_reg[48]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[48]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[56]_i_1 
       (.CI(\frame_128_255_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_128_255_transed_reg[56]_i_1_CO_UNCONNECTED [7],\frame_128_255_transed_reg[56]_i_1_n_1 ,\frame_128_255_transed_reg[56]_i_1_n_2 ,\frame_128_255_transed_reg[56]_i_1_n_3 ,\frame_128_255_transed_reg[56]_i_1_n_4 ,\frame_128_255_transed_reg[56]_i_1_n_5 ,\frame_128_255_transed_reg[56]_i_1_n_6 ,\frame_128_255_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[56]_i_1_n_8 ,\frame_128_255_transed_reg[56]_i_1_n_9 ,\frame_128_255_transed_reg[56]_i_1_n_10 ,\frame_128_255_transed_reg[56]_i_1_n_11 ,\frame_128_255_transed_reg[56]_i_1_n_12 ,\frame_128_255_transed_reg[56]_i_1_n_13 ,\frame_128_255_transed_reg[56]_i_1_n_14 ,\frame_128_255_transed_reg[56]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_13 ),
        .Q(frame_128_255_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_12 ),
        .Q(frame_128_255_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_11 ),
        .Q(frame_128_255_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_10 ),
        .Q(frame_128_255_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[56]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_9 ),
        .Q(frame_128_255_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[0]_i_1_n_8 ),
        .Q(frame_128_255_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_15 ),
        .Q(frame_128_255_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_128_255_transed_reg[8]_i_1 
       (.CI(\frame_128_255_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_128_255_transed_reg[8]_i_1_n_0 ,\frame_128_255_transed_reg[8]_i_1_n_1 ,\frame_128_255_transed_reg[8]_i_1_n_2 ,\frame_128_255_transed_reg[8]_i_1_n_3 ,\frame_128_255_transed_reg[8]_i_1_n_4 ,\frame_128_255_transed_reg[8]_i_1_n_5 ,\frame_128_255_transed_reg[8]_i_1_n_6 ,\frame_128_255_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_128_255_transed_reg[8]_i_1_n_8 ,\frame_128_255_transed_reg[8]_i_1_n_9 ,\frame_128_255_transed_reg[8]_i_1_n_10 ,\frame_128_255_transed_reg[8]_i_1_n_11 ,\frame_128_255_transed_reg[8]_i_1_n_12 ,\frame_128_255_transed_reg[8]_i_1_n_13 ,\frame_128_255_transed_reg[8]_i_1_n_14 ,\frame_128_255_transed_reg[8]_i_1_n_15 }),
        .S(frame_128_255_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_128_255_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_128_255_transed_reg[8]_i_1_n_14 ),
        .Q(frame_128_255_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_256_511_good[0]_i_2 
       (.I0(frame_256_511_good_reg[0]),
        .O(\frame_256_511_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[0]_i_1_n_0 ,\frame_256_511_good_reg[0]_i_1_n_1 ,\frame_256_511_good_reg[0]_i_1_n_2 ,\frame_256_511_good_reg[0]_i_1_n_3 ,\frame_256_511_good_reg[0]_i_1_n_4 ,\frame_256_511_good_reg[0]_i_1_n_5 ,\frame_256_511_good_reg[0]_i_1_n_6 ,\frame_256_511_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_256_511_good_reg[0]_i_1_n_8 ,\frame_256_511_good_reg[0]_i_1_n_9 ,\frame_256_511_good_reg[0]_i_1_n_10 ,\frame_256_511_good_reg[0]_i_1_n_11 ,\frame_256_511_good_reg[0]_i_1_n_12 ,\frame_256_511_good_reg[0]_i_1_n_13 ,\frame_256_511_good_reg[0]_i_1_n_14 ,\frame_256_511_good_reg[0]_i_1_n_15 }),
        .S({frame_256_511_good_reg[7:1],\frame_256_511_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[16]_i_1 
       (.CI(\frame_256_511_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[16]_i_1_n_0 ,\frame_256_511_good_reg[16]_i_1_n_1 ,\frame_256_511_good_reg[16]_i_1_n_2 ,\frame_256_511_good_reg[16]_i_1_n_3 ,\frame_256_511_good_reg[16]_i_1_n_4 ,\frame_256_511_good_reg[16]_i_1_n_5 ,\frame_256_511_good_reg[16]_i_1_n_6 ,\frame_256_511_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[16]_i_1_n_8 ,\frame_256_511_good_reg[16]_i_1_n_9 ,\frame_256_511_good_reg[16]_i_1_n_10 ,\frame_256_511_good_reg[16]_i_1_n_11 ,\frame_256_511_good_reg[16]_i_1_n_12 ,\frame_256_511_good_reg[16]_i_1_n_13 ,\frame_256_511_good_reg[16]_i_1_n_14 ,\frame_256_511_good_reg[16]_i_1_n_15 }),
        .S(frame_256_511_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[16]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[24]_i_1 
       (.CI(\frame_256_511_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[24]_i_1_n_0 ,\frame_256_511_good_reg[24]_i_1_n_1 ,\frame_256_511_good_reg[24]_i_1_n_2 ,\frame_256_511_good_reg[24]_i_1_n_3 ,\frame_256_511_good_reg[24]_i_1_n_4 ,\frame_256_511_good_reg[24]_i_1_n_5 ,\frame_256_511_good_reg[24]_i_1_n_6 ,\frame_256_511_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[24]_i_1_n_8 ,\frame_256_511_good_reg[24]_i_1_n_9 ,\frame_256_511_good_reg[24]_i_1_n_10 ,\frame_256_511_good_reg[24]_i_1_n_11 ,\frame_256_511_good_reg[24]_i_1_n_12 ,\frame_256_511_good_reg[24]_i_1_n_13 ,\frame_256_511_good_reg[24]_i_1_n_14 ,\frame_256_511_good_reg[24]_i_1_n_15 }),
        .S(frame_256_511_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[24]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[32]_i_1 
       (.CI(\frame_256_511_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[32]_i_1_n_0 ,\frame_256_511_good_reg[32]_i_1_n_1 ,\frame_256_511_good_reg[32]_i_1_n_2 ,\frame_256_511_good_reg[32]_i_1_n_3 ,\frame_256_511_good_reg[32]_i_1_n_4 ,\frame_256_511_good_reg[32]_i_1_n_5 ,\frame_256_511_good_reg[32]_i_1_n_6 ,\frame_256_511_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[32]_i_1_n_8 ,\frame_256_511_good_reg[32]_i_1_n_9 ,\frame_256_511_good_reg[32]_i_1_n_10 ,\frame_256_511_good_reg[32]_i_1_n_11 ,\frame_256_511_good_reg[32]_i_1_n_12 ,\frame_256_511_good_reg[32]_i_1_n_13 ,\frame_256_511_good_reg[32]_i_1_n_14 ,\frame_256_511_good_reg[32]_i_1_n_15 }),
        .S(frame_256_511_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[32]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[40]_i_1 
       (.CI(\frame_256_511_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[40]_i_1_n_0 ,\frame_256_511_good_reg[40]_i_1_n_1 ,\frame_256_511_good_reg[40]_i_1_n_2 ,\frame_256_511_good_reg[40]_i_1_n_3 ,\frame_256_511_good_reg[40]_i_1_n_4 ,\frame_256_511_good_reg[40]_i_1_n_5 ,\frame_256_511_good_reg[40]_i_1_n_6 ,\frame_256_511_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[40]_i_1_n_8 ,\frame_256_511_good_reg[40]_i_1_n_9 ,\frame_256_511_good_reg[40]_i_1_n_10 ,\frame_256_511_good_reg[40]_i_1_n_11 ,\frame_256_511_good_reg[40]_i_1_n_12 ,\frame_256_511_good_reg[40]_i_1_n_13 ,\frame_256_511_good_reg[40]_i_1_n_14 ,\frame_256_511_good_reg[40]_i_1_n_15 }),
        .S(frame_256_511_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[40]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[48]_i_1 
       (.CI(\frame_256_511_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[48]_i_1_n_0 ,\frame_256_511_good_reg[48]_i_1_n_1 ,\frame_256_511_good_reg[48]_i_1_n_2 ,\frame_256_511_good_reg[48]_i_1_n_3 ,\frame_256_511_good_reg[48]_i_1_n_4 ,\frame_256_511_good_reg[48]_i_1_n_5 ,\frame_256_511_good_reg[48]_i_1_n_6 ,\frame_256_511_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[48]_i_1_n_8 ,\frame_256_511_good_reg[48]_i_1_n_9 ,\frame_256_511_good_reg[48]_i_1_n_10 ,\frame_256_511_good_reg[48]_i_1_n_11 ,\frame_256_511_good_reg[48]_i_1_n_12 ,\frame_256_511_good_reg[48]_i_1_n_13 ,\frame_256_511_good_reg[48]_i_1_n_14 ,\frame_256_511_good_reg[48]_i_1_n_15 }),
        .S(frame_256_511_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[48]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[56]_i_1 
       (.CI(\frame_256_511_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_256_511_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_256_511_good_reg[56]_i_1_n_1 ,\frame_256_511_good_reg[56]_i_1_n_2 ,\frame_256_511_good_reg[56]_i_1_n_3 ,\frame_256_511_good_reg[56]_i_1_n_4 ,\frame_256_511_good_reg[56]_i_1_n_5 ,\frame_256_511_good_reg[56]_i_1_n_6 ,\frame_256_511_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[56]_i_1_n_8 ,\frame_256_511_good_reg[56]_i_1_n_9 ,\frame_256_511_good_reg[56]_i_1_n_10 ,\frame_256_511_good_reg[56]_i_1_n_11 ,\frame_256_511_good_reg[56]_i_1_n_12 ,\frame_256_511_good_reg[56]_i_1_n_13 ,\frame_256_511_good_reg[56]_i_1_n_14 ,\frame_256_511_good_reg[56]_i_1_n_15 }),
        .S(frame_256_511_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_13 ),
        .Q(frame_256_511_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_12 ),
        .Q(frame_256_511_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_11 ),
        .Q(frame_256_511_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_10 ),
        .Q(frame_256_511_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[56]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_9 ),
        .Q(frame_256_511_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[0]_i_1_n_8 ),
        .Q(frame_256_511_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_15 ),
        .Q(frame_256_511_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_good_reg[8]_i_1 
       (.CI(\frame_256_511_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_good_reg[8]_i_1_n_0 ,\frame_256_511_good_reg[8]_i_1_n_1 ,\frame_256_511_good_reg[8]_i_1_n_2 ,\frame_256_511_good_reg[8]_i_1_n_3 ,\frame_256_511_good_reg[8]_i_1_n_4 ,\frame_256_511_good_reg[8]_i_1_n_5 ,\frame_256_511_good_reg[8]_i_1_n_6 ,\frame_256_511_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_good_reg[8]_i_1_n_8 ,\frame_256_511_good_reg[8]_i_1_n_9 ,\frame_256_511_good_reg[8]_i_1_n_10 ,\frame_256_511_good_reg[8]_i_1_n_11 ,\frame_256_511_good_reg[8]_i_1_n_12 ,\frame_256_511_good_reg[8]_i_1_n_13 ,\frame_256_511_good_reg[8]_i_1_n_14 ,\frame_256_511_good_reg[8]_i_1_n_15 }),
        .S(frame_256_511_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_256_511_good_reg[8]_i_1_n_14 ),
        .Q(frame_256_511_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_256_511_transed[0]_i_2 
       (.I0(frame_256_511_transed_reg[0]),
        .O(\frame_256_511_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[0]_i_1_n_0 ,\frame_256_511_transed_reg[0]_i_1_n_1 ,\frame_256_511_transed_reg[0]_i_1_n_2 ,\frame_256_511_transed_reg[0]_i_1_n_3 ,\frame_256_511_transed_reg[0]_i_1_n_4 ,\frame_256_511_transed_reg[0]_i_1_n_5 ,\frame_256_511_transed_reg[0]_i_1_n_6 ,\frame_256_511_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_256_511_transed_reg[0]_i_1_n_8 ,\frame_256_511_transed_reg[0]_i_1_n_9 ,\frame_256_511_transed_reg[0]_i_1_n_10 ,\frame_256_511_transed_reg[0]_i_1_n_11 ,\frame_256_511_transed_reg[0]_i_1_n_12 ,\frame_256_511_transed_reg[0]_i_1_n_13 ,\frame_256_511_transed_reg[0]_i_1_n_14 ,\frame_256_511_transed_reg[0]_i_1_n_15 }),
        .S({frame_256_511_transed_reg[7:1],\frame_256_511_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[16]_i_1 
       (.CI(\frame_256_511_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[16]_i_1_n_0 ,\frame_256_511_transed_reg[16]_i_1_n_1 ,\frame_256_511_transed_reg[16]_i_1_n_2 ,\frame_256_511_transed_reg[16]_i_1_n_3 ,\frame_256_511_transed_reg[16]_i_1_n_4 ,\frame_256_511_transed_reg[16]_i_1_n_5 ,\frame_256_511_transed_reg[16]_i_1_n_6 ,\frame_256_511_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[16]_i_1_n_8 ,\frame_256_511_transed_reg[16]_i_1_n_9 ,\frame_256_511_transed_reg[16]_i_1_n_10 ,\frame_256_511_transed_reg[16]_i_1_n_11 ,\frame_256_511_transed_reg[16]_i_1_n_12 ,\frame_256_511_transed_reg[16]_i_1_n_13 ,\frame_256_511_transed_reg[16]_i_1_n_14 ,\frame_256_511_transed_reg[16]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[16]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[24]_i_1 
       (.CI(\frame_256_511_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[24]_i_1_n_0 ,\frame_256_511_transed_reg[24]_i_1_n_1 ,\frame_256_511_transed_reg[24]_i_1_n_2 ,\frame_256_511_transed_reg[24]_i_1_n_3 ,\frame_256_511_transed_reg[24]_i_1_n_4 ,\frame_256_511_transed_reg[24]_i_1_n_5 ,\frame_256_511_transed_reg[24]_i_1_n_6 ,\frame_256_511_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[24]_i_1_n_8 ,\frame_256_511_transed_reg[24]_i_1_n_9 ,\frame_256_511_transed_reg[24]_i_1_n_10 ,\frame_256_511_transed_reg[24]_i_1_n_11 ,\frame_256_511_transed_reg[24]_i_1_n_12 ,\frame_256_511_transed_reg[24]_i_1_n_13 ,\frame_256_511_transed_reg[24]_i_1_n_14 ,\frame_256_511_transed_reg[24]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[24]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[32]_i_1 
       (.CI(\frame_256_511_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[32]_i_1_n_0 ,\frame_256_511_transed_reg[32]_i_1_n_1 ,\frame_256_511_transed_reg[32]_i_1_n_2 ,\frame_256_511_transed_reg[32]_i_1_n_3 ,\frame_256_511_transed_reg[32]_i_1_n_4 ,\frame_256_511_transed_reg[32]_i_1_n_5 ,\frame_256_511_transed_reg[32]_i_1_n_6 ,\frame_256_511_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[32]_i_1_n_8 ,\frame_256_511_transed_reg[32]_i_1_n_9 ,\frame_256_511_transed_reg[32]_i_1_n_10 ,\frame_256_511_transed_reg[32]_i_1_n_11 ,\frame_256_511_transed_reg[32]_i_1_n_12 ,\frame_256_511_transed_reg[32]_i_1_n_13 ,\frame_256_511_transed_reg[32]_i_1_n_14 ,\frame_256_511_transed_reg[32]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[32]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[40]_i_1 
       (.CI(\frame_256_511_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[40]_i_1_n_0 ,\frame_256_511_transed_reg[40]_i_1_n_1 ,\frame_256_511_transed_reg[40]_i_1_n_2 ,\frame_256_511_transed_reg[40]_i_1_n_3 ,\frame_256_511_transed_reg[40]_i_1_n_4 ,\frame_256_511_transed_reg[40]_i_1_n_5 ,\frame_256_511_transed_reg[40]_i_1_n_6 ,\frame_256_511_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[40]_i_1_n_8 ,\frame_256_511_transed_reg[40]_i_1_n_9 ,\frame_256_511_transed_reg[40]_i_1_n_10 ,\frame_256_511_transed_reg[40]_i_1_n_11 ,\frame_256_511_transed_reg[40]_i_1_n_12 ,\frame_256_511_transed_reg[40]_i_1_n_13 ,\frame_256_511_transed_reg[40]_i_1_n_14 ,\frame_256_511_transed_reg[40]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[40]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[48]_i_1 
       (.CI(\frame_256_511_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[48]_i_1_n_0 ,\frame_256_511_transed_reg[48]_i_1_n_1 ,\frame_256_511_transed_reg[48]_i_1_n_2 ,\frame_256_511_transed_reg[48]_i_1_n_3 ,\frame_256_511_transed_reg[48]_i_1_n_4 ,\frame_256_511_transed_reg[48]_i_1_n_5 ,\frame_256_511_transed_reg[48]_i_1_n_6 ,\frame_256_511_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[48]_i_1_n_8 ,\frame_256_511_transed_reg[48]_i_1_n_9 ,\frame_256_511_transed_reg[48]_i_1_n_10 ,\frame_256_511_transed_reg[48]_i_1_n_11 ,\frame_256_511_transed_reg[48]_i_1_n_12 ,\frame_256_511_transed_reg[48]_i_1_n_13 ,\frame_256_511_transed_reg[48]_i_1_n_14 ,\frame_256_511_transed_reg[48]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[48]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[56]_i_1 
       (.CI(\frame_256_511_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_256_511_transed_reg[56]_i_1_CO_UNCONNECTED [7],\frame_256_511_transed_reg[56]_i_1_n_1 ,\frame_256_511_transed_reg[56]_i_1_n_2 ,\frame_256_511_transed_reg[56]_i_1_n_3 ,\frame_256_511_transed_reg[56]_i_1_n_4 ,\frame_256_511_transed_reg[56]_i_1_n_5 ,\frame_256_511_transed_reg[56]_i_1_n_6 ,\frame_256_511_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[56]_i_1_n_8 ,\frame_256_511_transed_reg[56]_i_1_n_9 ,\frame_256_511_transed_reg[56]_i_1_n_10 ,\frame_256_511_transed_reg[56]_i_1_n_11 ,\frame_256_511_transed_reg[56]_i_1_n_12 ,\frame_256_511_transed_reg[56]_i_1_n_13 ,\frame_256_511_transed_reg[56]_i_1_n_14 ,\frame_256_511_transed_reg[56]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_13 ),
        .Q(frame_256_511_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_12 ),
        .Q(frame_256_511_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_11 ),
        .Q(frame_256_511_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_10 ),
        .Q(frame_256_511_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[56]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_9 ),
        .Q(frame_256_511_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[0]_i_1_n_8 ),
        .Q(frame_256_511_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_15 ),
        .Q(frame_256_511_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_256_511_transed_reg[8]_i_1 
       (.CI(\frame_256_511_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_256_511_transed_reg[8]_i_1_n_0 ,\frame_256_511_transed_reg[8]_i_1_n_1 ,\frame_256_511_transed_reg[8]_i_1_n_2 ,\frame_256_511_transed_reg[8]_i_1_n_3 ,\frame_256_511_transed_reg[8]_i_1_n_4 ,\frame_256_511_transed_reg[8]_i_1_n_5 ,\frame_256_511_transed_reg[8]_i_1_n_6 ,\frame_256_511_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_256_511_transed_reg[8]_i_1_n_8 ,\frame_256_511_transed_reg[8]_i_1_n_9 ,\frame_256_511_transed_reg[8]_i_1_n_10 ,\frame_256_511_transed_reg[8]_i_1_n_11 ,\frame_256_511_transed_reg[8]_i_1_n_12 ,\frame_256_511_transed_reg[8]_i_1_n_13 ,\frame_256_511_transed_reg[8]_i_1_n_14 ,\frame_256_511_transed_reg[8]_i_1_n_15 }),
        .S(frame_256_511_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_256_511_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[9]),
        .CLR(rst_i),
        .D(\frame_256_511_transed_reg[8]_i_1_n_14 ),
        .Q(frame_256_511_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_512_1023_good[0]_i_2 
       (.I0(frame_512_1023_good_reg[0]),
        .O(\frame_512_1023_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[0]_i_1_n_0 ,\frame_512_1023_good_reg[0]_i_1_n_1 ,\frame_512_1023_good_reg[0]_i_1_n_2 ,\frame_512_1023_good_reg[0]_i_1_n_3 ,\frame_512_1023_good_reg[0]_i_1_n_4 ,\frame_512_1023_good_reg[0]_i_1_n_5 ,\frame_512_1023_good_reg[0]_i_1_n_6 ,\frame_512_1023_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_512_1023_good_reg[0]_i_1_n_8 ,\frame_512_1023_good_reg[0]_i_1_n_9 ,\frame_512_1023_good_reg[0]_i_1_n_10 ,\frame_512_1023_good_reg[0]_i_1_n_11 ,\frame_512_1023_good_reg[0]_i_1_n_12 ,\frame_512_1023_good_reg[0]_i_1_n_13 ,\frame_512_1023_good_reg[0]_i_1_n_14 ,\frame_512_1023_good_reg[0]_i_1_n_15 }),
        .S({frame_512_1023_good_reg[7:1],\frame_512_1023_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[16]_i_1 
       (.CI(\frame_512_1023_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[16]_i_1_n_0 ,\frame_512_1023_good_reg[16]_i_1_n_1 ,\frame_512_1023_good_reg[16]_i_1_n_2 ,\frame_512_1023_good_reg[16]_i_1_n_3 ,\frame_512_1023_good_reg[16]_i_1_n_4 ,\frame_512_1023_good_reg[16]_i_1_n_5 ,\frame_512_1023_good_reg[16]_i_1_n_6 ,\frame_512_1023_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[16]_i_1_n_8 ,\frame_512_1023_good_reg[16]_i_1_n_9 ,\frame_512_1023_good_reg[16]_i_1_n_10 ,\frame_512_1023_good_reg[16]_i_1_n_11 ,\frame_512_1023_good_reg[16]_i_1_n_12 ,\frame_512_1023_good_reg[16]_i_1_n_13 ,\frame_512_1023_good_reg[16]_i_1_n_14 ,\frame_512_1023_good_reg[16]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[16]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[24]_i_1 
       (.CI(\frame_512_1023_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[24]_i_1_n_0 ,\frame_512_1023_good_reg[24]_i_1_n_1 ,\frame_512_1023_good_reg[24]_i_1_n_2 ,\frame_512_1023_good_reg[24]_i_1_n_3 ,\frame_512_1023_good_reg[24]_i_1_n_4 ,\frame_512_1023_good_reg[24]_i_1_n_5 ,\frame_512_1023_good_reg[24]_i_1_n_6 ,\frame_512_1023_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[24]_i_1_n_8 ,\frame_512_1023_good_reg[24]_i_1_n_9 ,\frame_512_1023_good_reg[24]_i_1_n_10 ,\frame_512_1023_good_reg[24]_i_1_n_11 ,\frame_512_1023_good_reg[24]_i_1_n_12 ,\frame_512_1023_good_reg[24]_i_1_n_13 ,\frame_512_1023_good_reg[24]_i_1_n_14 ,\frame_512_1023_good_reg[24]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[24]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[32]_i_1 
       (.CI(\frame_512_1023_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[32]_i_1_n_0 ,\frame_512_1023_good_reg[32]_i_1_n_1 ,\frame_512_1023_good_reg[32]_i_1_n_2 ,\frame_512_1023_good_reg[32]_i_1_n_3 ,\frame_512_1023_good_reg[32]_i_1_n_4 ,\frame_512_1023_good_reg[32]_i_1_n_5 ,\frame_512_1023_good_reg[32]_i_1_n_6 ,\frame_512_1023_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[32]_i_1_n_8 ,\frame_512_1023_good_reg[32]_i_1_n_9 ,\frame_512_1023_good_reg[32]_i_1_n_10 ,\frame_512_1023_good_reg[32]_i_1_n_11 ,\frame_512_1023_good_reg[32]_i_1_n_12 ,\frame_512_1023_good_reg[32]_i_1_n_13 ,\frame_512_1023_good_reg[32]_i_1_n_14 ,\frame_512_1023_good_reg[32]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[32]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[40]_i_1 
       (.CI(\frame_512_1023_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[40]_i_1_n_0 ,\frame_512_1023_good_reg[40]_i_1_n_1 ,\frame_512_1023_good_reg[40]_i_1_n_2 ,\frame_512_1023_good_reg[40]_i_1_n_3 ,\frame_512_1023_good_reg[40]_i_1_n_4 ,\frame_512_1023_good_reg[40]_i_1_n_5 ,\frame_512_1023_good_reg[40]_i_1_n_6 ,\frame_512_1023_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[40]_i_1_n_8 ,\frame_512_1023_good_reg[40]_i_1_n_9 ,\frame_512_1023_good_reg[40]_i_1_n_10 ,\frame_512_1023_good_reg[40]_i_1_n_11 ,\frame_512_1023_good_reg[40]_i_1_n_12 ,\frame_512_1023_good_reg[40]_i_1_n_13 ,\frame_512_1023_good_reg[40]_i_1_n_14 ,\frame_512_1023_good_reg[40]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[40]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[48]_i_1 
       (.CI(\frame_512_1023_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[48]_i_1_n_0 ,\frame_512_1023_good_reg[48]_i_1_n_1 ,\frame_512_1023_good_reg[48]_i_1_n_2 ,\frame_512_1023_good_reg[48]_i_1_n_3 ,\frame_512_1023_good_reg[48]_i_1_n_4 ,\frame_512_1023_good_reg[48]_i_1_n_5 ,\frame_512_1023_good_reg[48]_i_1_n_6 ,\frame_512_1023_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[48]_i_1_n_8 ,\frame_512_1023_good_reg[48]_i_1_n_9 ,\frame_512_1023_good_reg[48]_i_1_n_10 ,\frame_512_1023_good_reg[48]_i_1_n_11 ,\frame_512_1023_good_reg[48]_i_1_n_12 ,\frame_512_1023_good_reg[48]_i_1_n_13 ,\frame_512_1023_good_reg[48]_i_1_n_14 ,\frame_512_1023_good_reg[48]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[48]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[56]_i_1 
       (.CI(\frame_512_1023_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_512_1023_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_512_1023_good_reg[56]_i_1_n_1 ,\frame_512_1023_good_reg[56]_i_1_n_2 ,\frame_512_1023_good_reg[56]_i_1_n_3 ,\frame_512_1023_good_reg[56]_i_1_n_4 ,\frame_512_1023_good_reg[56]_i_1_n_5 ,\frame_512_1023_good_reg[56]_i_1_n_6 ,\frame_512_1023_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[56]_i_1_n_8 ,\frame_512_1023_good_reg[56]_i_1_n_9 ,\frame_512_1023_good_reg[56]_i_1_n_10 ,\frame_512_1023_good_reg[56]_i_1_n_11 ,\frame_512_1023_good_reg[56]_i_1_n_12 ,\frame_512_1023_good_reg[56]_i_1_n_13 ,\frame_512_1023_good_reg[56]_i_1_n_14 ,\frame_512_1023_good_reg[56]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_13 ),
        .Q(frame_512_1023_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_12 ),
        .Q(frame_512_1023_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_11 ),
        .Q(frame_512_1023_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_10 ),
        .Q(frame_512_1023_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[56]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_9 ),
        .Q(frame_512_1023_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[0]_i_1_n_8 ),
        .Q(frame_512_1023_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_15 ),
        .Q(frame_512_1023_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_good_reg[8]_i_1 
       (.CI(\frame_512_1023_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_good_reg[8]_i_1_n_0 ,\frame_512_1023_good_reg[8]_i_1_n_1 ,\frame_512_1023_good_reg[8]_i_1_n_2 ,\frame_512_1023_good_reg[8]_i_1_n_3 ,\frame_512_1023_good_reg[8]_i_1_n_4 ,\frame_512_1023_good_reg[8]_i_1_n_5 ,\frame_512_1023_good_reg[8]_i_1_n_6 ,\frame_512_1023_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_good_reg[8]_i_1_n_8 ,\frame_512_1023_good_reg[8]_i_1_n_9 ,\frame_512_1023_good_reg[8]_i_1_n_10 ,\frame_512_1023_good_reg[8]_i_1_n_11 ,\frame_512_1023_good_reg[8]_i_1_n_12 ,\frame_512_1023_good_reg[8]_i_1_n_13 ,\frame_512_1023_good_reg[8]_i_1_n_14 ,\frame_512_1023_good_reg[8]_i_1_n_15 }),
        .S(frame_512_1023_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[8]),
        .CLR(rst_i),
        .D(\frame_512_1023_good_reg[8]_i_1_n_14 ),
        .Q(frame_512_1023_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_512_1023_transed[0]_i_2 
       (.I0(frame_512_1023_transed_reg[0]),
        .O(\frame_512_1023_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[0]_i_1_n_0 ,\frame_512_1023_transed_reg[0]_i_1_n_1 ,\frame_512_1023_transed_reg[0]_i_1_n_2 ,\frame_512_1023_transed_reg[0]_i_1_n_3 ,\frame_512_1023_transed_reg[0]_i_1_n_4 ,\frame_512_1023_transed_reg[0]_i_1_n_5 ,\frame_512_1023_transed_reg[0]_i_1_n_6 ,\frame_512_1023_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_512_1023_transed_reg[0]_i_1_n_8 ,\frame_512_1023_transed_reg[0]_i_1_n_9 ,\frame_512_1023_transed_reg[0]_i_1_n_10 ,\frame_512_1023_transed_reg[0]_i_1_n_11 ,\frame_512_1023_transed_reg[0]_i_1_n_12 ,\frame_512_1023_transed_reg[0]_i_1_n_13 ,\frame_512_1023_transed_reg[0]_i_1_n_14 ,\frame_512_1023_transed_reg[0]_i_1_n_15 }),
        .S({frame_512_1023_transed_reg[7:1],\frame_512_1023_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[16]_i_1 
       (.CI(\frame_512_1023_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[16]_i_1_n_0 ,\frame_512_1023_transed_reg[16]_i_1_n_1 ,\frame_512_1023_transed_reg[16]_i_1_n_2 ,\frame_512_1023_transed_reg[16]_i_1_n_3 ,\frame_512_1023_transed_reg[16]_i_1_n_4 ,\frame_512_1023_transed_reg[16]_i_1_n_5 ,\frame_512_1023_transed_reg[16]_i_1_n_6 ,\frame_512_1023_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[16]_i_1_n_8 ,\frame_512_1023_transed_reg[16]_i_1_n_9 ,\frame_512_1023_transed_reg[16]_i_1_n_10 ,\frame_512_1023_transed_reg[16]_i_1_n_11 ,\frame_512_1023_transed_reg[16]_i_1_n_12 ,\frame_512_1023_transed_reg[16]_i_1_n_13 ,\frame_512_1023_transed_reg[16]_i_1_n_14 ,\frame_512_1023_transed_reg[16]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[16]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[24]_i_1 
       (.CI(\frame_512_1023_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[24]_i_1_n_0 ,\frame_512_1023_transed_reg[24]_i_1_n_1 ,\frame_512_1023_transed_reg[24]_i_1_n_2 ,\frame_512_1023_transed_reg[24]_i_1_n_3 ,\frame_512_1023_transed_reg[24]_i_1_n_4 ,\frame_512_1023_transed_reg[24]_i_1_n_5 ,\frame_512_1023_transed_reg[24]_i_1_n_6 ,\frame_512_1023_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[24]_i_1_n_8 ,\frame_512_1023_transed_reg[24]_i_1_n_9 ,\frame_512_1023_transed_reg[24]_i_1_n_10 ,\frame_512_1023_transed_reg[24]_i_1_n_11 ,\frame_512_1023_transed_reg[24]_i_1_n_12 ,\frame_512_1023_transed_reg[24]_i_1_n_13 ,\frame_512_1023_transed_reg[24]_i_1_n_14 ,\frame_512_1023_transed_reg[24]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[24]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[32]_i_1 
       (.CI(\frame_512_1023_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[32]_i_1_n_0 ,\frame_512_1023_transed_reg[32]_i_1_n_1 ,\frame_512_1023_transed_reg[32]_i_1_n_2 ,\frame_512_1023_transed_reg[32]_i_1_n_3 ,\frame_512_1023_transed_reg[32]_i_1_n_4 ,\frame_512_1023_transed_reg[32]_i_1_n_5 ,\frame_512_1023_transed_reg[32]_i_1_n_6 ,\frame_512_1023_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[32]_i_1_n_8 ,\frame_512_1023_transed_reg[32]_i_1_n_9 ,\frame_512_1023_transed_reg[32]_i_1_n_10 ,\frame_512_1023_transed_reg[32]_i_1_n_11 ,\frame_512_1023_transed_reg[32]_i_1_n_12 ,\frame_512_1023_transed_reg[32]_i_1_n_13 ,\frame_512_1023_transed_reg[32]_i_1_n_14 ,\frame_512_1023_transed_reg[32]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[32]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[40]_i_1 
       (.CI(\frame_512_1023_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[40]_i_1_n_0 ,\frame_512_1023_transed_reg[40]_i_1_n_1 ,\frame_512_1023_transed_reg[40]_i_1_n_2 ,\frame_512_1023_transed_reg[40]_i_1_n_3 ,\frame_512_1023_transed_reg[40]_i_1_n_4 ,\frame_512_1023_transed_reg[40]_i_1_n_5 ,\frame_512_1023_transed_reg[40]_i_1_n_6 ,\frame_512_1023_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[40]_i_1_n_8 ,\frame_512_1023_transed_reg[40]_i_1_n_9 ,\frame_512_1023_transed_reg[40]_i_1_n_10 ,\frame_512_1023_transed_reg[40]_i_1_n_11 ,\frame_512_1023_transed_reg[40]_i_1_n_12 ,\frame_512_1023_transed_reg[40]_i_1_n_13 ,\frame_512_1023_transed_reg[40]_i_1_n_14 ,\frame_512_1023_transed_reg[40]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[40]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[48]_i_1 
       (.CI(\frame_512_1023_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[48]_i_1_n_0 ,\frame_512_1023_transed_reg[48]_i_1_n_1 ,\frame_512_1023_transed_reg[48]_i_1_n_2 ,\frame_512_1023_transed_reg[48]_i_1_n_3 ,\frame_512_1023_transed_reg[48]_i_1_n_4 ,\frame_512_1023_transed_reg[48]_i_1_n_5 ,\frame_512_1023_transed_reg[48]_i_1_n_6 ,\frame_512_1023_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[48]_i_1_n_8 ,\frame_512_1023_transed_reg[48]_i_1_n_9 ,\frame_512_1023_transed_reg[48]_i_1_n_10 ,\frame_512_1023_transed_reg[48]_i_1_n_11 ,\frame_512_1023_transed_reg[48]_i_1_n_12 ,\frame_512_1023_transed_reg[48]_i_1_n_13 ,\frame_512_1023_transed_reg[48]_i_1_n_14 ,\frame_512_1023_transed_reg[48]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[48]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[56]_i_1 
       (.CI(\frame_512_1023_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_512_1023_transed_reg[56]_i_1_CO_UNCONNECTED [7],\frame_512_1023_transed_reg[56]_i_1_n_1 ,\frame_512_1023_transed_reg[56]_i_1_n_2 ,\frame_512_1023_transed_reg[56]_i_1_n_3 ,\frame_512_1023_transed_reg[56]_i_1_n_4 ,\frame_512_1023_transed_reg[56]_i_1_n_5 ,\frame_512_1023_transed_reg[56]_i_1_n_6 ,\frame_512_1023_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[56]_i_1_n_8 ,\frame_512_1023_transed_reg[56]_i_1_n_9 ,\frame_512_1023_transed_reg[56]_i_1_n_10 ,\frame_512_1023_transed_reg[56]_i_1_n_11 ,\frame_512_1023_transed_reg[56]_i_1_n_12 ,\frame_512_1023_transed_reg[56]_i_1_n_13 ,\frame_512_1023_transed_reg[56]_i_1_n_14 ,\frame_512_1023_transed_reg[56]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_13 ),
        .Q(frame_512_1023_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_12 ),
        .Q(frame_512_1023_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_11 ),
        .Q(frame_512_1023_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_10 ),
        .Q(frame_512_1023_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[56]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_9 ),
        .Q(frame_512_1023_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[0]_i_1_n_8 ),
        .Q(frame_512_1023_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_15 ),
        .Q(frame_512_1023_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_512_1023_transed_reg[8]_i_1 
       (.CI(\frame_512_1023_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_512_1023_transed_reg[8]_i_1_n_0 ,\frame_512_1023_transed_reg[8]_i_1_n_1 ,\frame_512_1023_transed_reg[8]_i_1_n_2 ,\frame_512_1023_transed_reg[8]_i_1_n_3 ,\frame_512_1023_transed_reg[8]_i_1_n_4 ,\frame_512_1023_transed_reg[8]_i_1_n_5 ,\frame_512_1023_transed_reg[8]_i_1_n_6 ,\frame_512_1023_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_512_1023_transed_reg[8]_i_1_n_8 ,\frame_512_1023_transed_reg[8]_i_1_n_9 ,\frame_512_1023_transed_reg[8]_i_1_n_10 ,\frame_512_1023_transed_reg[8]_i_1_n_11 ,\frame_512_1023_transed_reg[8]_i_1_n_12 ,\frame_512_1023_transed_reg[8]_i_1_n_13 ,\frame_512_1023_transed_reg[8]_i_1_n_14 ,\frame_512_1023_transed_reg[8]_i_1_n_15 }),
        .S(frame_512_1023_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_512_1023_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[10]),
        .CLR(rst_i),
        .D(\frame_512_1023_transed_reg[8]_i_1_n_14 ),
        .Q(frame_512_1023_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_64_good[0]_i_2 
       (.I0(frame_64_good_reg[0]),
        .O(\frame_64_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_15 ),
        .Q(frame_64_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[0]_i_1_n_0 ,\frame_64_good_reg[0]_i_1_n_1 ,\frame_64_good_reg[0]_i_1_n_2 ,\frame_64_good_reg[0]_i_1_n_3 ,\frame_64_good_reg[0]_i_1_n_4 ,\frame_64_good_reg[0]_i_1_n_5 ,\frame_64_good_reg[0]_i_1_n_6 ,\frame_64_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_64_good_reg[0]_i_1_n_8 ,\frame_64_good_reg[0]_i_1_n_9 ,\frame_64_good_reg[0]_i_1_n_10 ,\frame_64_good_reg[0]_i_1_n_11 ,\frame_64_good_reg[0]_i_1_n_12 ,\frame_64_good_reg[0]_i_1_n_13 ,\frame_64_good_reg[0]_i_1_n_14 ,\frame_64_good_reg[0]_i_1_n_15 }),
        .S({frame_64_good_reg[7:1],\frame_64_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_13 ),
        .Q(frame_64_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_12 ),
        .Q(frame_64_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_11 ),
        .Q(frame_64_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_10 ),
        .Q(frame_64_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_9 ),
        .Q(frame_64_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_8 ),
        .Q(frame_64_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_15 ),
        .Q(frame_64_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[16]_i_1 
       (.CI(\frame_64_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[16]_i_1_n_0 ,\frame_64_good_reg[16]_i_1_n_1 ,\frame_64_good_reg[16]_i_1_n_2 ,\frame_64_good_reg[16]_i_1_n_3 ,\frame_64_good_reg[16]_i_1_n_4 ,\frame_64_good_reg[16]_i_1_n_5 ,\frame_64_good_reg[16]_i_1_n_6 ,\frame_64_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[16]_i_1_n_8 ,\frame_64_good_reg[16]_i_1_n_9 ,\frame_64_good_reg[16]_i_1_n_10 ,\frame_64_good_reg[16]_i_1_n_11 ,\frame_64_good_reg[16]_i_1_n_12 ,\frame_64_good_reg[16]_i_1_n_13 ,\frame_64_good_reg[16]_i_1_n_14 ,\frame_64_good_reg[16]_i_1_n_15 }),
        .S(frame_64_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_14 ),
        .Q(frame_64_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_13 ),
        .Q(frame_64_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_12 ),
        .Q(frame_64_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_14 ),
        .Q(frame_64_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_11 ),
        .Q(frame_64_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_10 ),
        .Q(frame_64_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_9 ),
        .Q(frame_64_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[16]_i_1_n_8 ),
        .Q(frame_64_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_15 ),
        .Q(frame_64_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[24]_i_1 
       (.CI(\frame_64_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[24]_i_1_n_0 ,\frame_64_good_reg[24]_i_1_n_1 ,\frame_64_good_reg[24]_i_1_n_2 ,\frame_64_good_reg[24]_i_1_n_3 ,\frame_64_good_reg[24]_i_1_n_4 ,\frame_64_good_reg[24]_i_1_n_5 ,\frame_64_good_reg[24]_i_1_n_6 ,\frame_64_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[24]_i_1_n_8 ,\frame_64_good_reg[24]_i_1_n_9 ,\frame_64_good_reg[24]_i_1_n_10 ,\frame_64_good_reg[24]_i_1_n_11 ,\frame_64_good_reg[24]_i_1_n_12 ,\frame_64_good_reg[24]_i_1_n_13 ,\frame_64_good_reg[24]_i_1_n_14 ,\frame_64_good_reg[24]_i_1_n_15 }),
        .S(frame_64_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_14 ),
        .Q(frame_64_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_13 ),
        .Q(frame_64_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_12 ),
        .Q(frame_64_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_11 ),
        .Q(frame_64_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_10 ),
        .Q(frame_64_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_13 ),
        .Q(frame_64_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_9 ),
        .Q(frame_64_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[24]_i_1_n_8 ),
        .Q(frame_64_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_15 ),
        .Q(frame_64_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[32]_i_1 
       (.CI(\frame_64_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[32]_i_1_n_0 ,\frame_64_good_reg[32]_i_1_n_1 ,\frame_64_good_reg[32]_i_1_n_2 ,\frame_64_good_reg[32]_i_1_n_3 ,\frame_64_good_reg[32]_i_1_n_4 ,\frame_64_good_reg[32]_i_1_n_5 ,\frame_64_good_reg[32]_i_1_n_6 ,\frame_64_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[32]_i_1_n_8 ,\frame_64_good_reg[32]_i_1_n_9 ,\frame_64_good_reg[32]_i_1_n_10 ,\frame_64_good_reg[32]_i_1_n_11 ,\frame_64_good_reg[32]_i_1_n_12 ,\frame_64_good_reg[32]_i_1_n_13 ,\frame_64_good_reg[32]_i_1_n_14 ,\frame_64_good_reg[32]_i_1_n_15 }),
        .S(frame_64_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_14 ),
        .Q(frame_64_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_13 ),
        .Q(frame_64_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_12 ),
        .Q(frame_64_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_11 ),
        .Q(frame_64_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_10 ),
        .Q(frame_64_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_9 ),
        .Q(frame_64_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[32]_i_1_n_8 ),
        .Q(frame_64_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_12 ),
        .Q(frame_64_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_15 ),
        .Q(frame_64_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[40]_i_1 
       (.CI(\frame_64_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[40]_i_1_n_0 ,\frame_64_good_reg[40]_i_1_n_1 ,\frame_64_good_reg[40]_i_1_n_2 ,\frame_64_good_reg[40]_i_1_n_3 ,\frame_64_good_reg[40]_i_1_n_4 ,\frame_64_good_reg[40]_i_1_n_5 ,\frame_64_good_reg[40]_i_1_n_6 ,\frame_64_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[40]_i_1_n_8 ,\frame_64_good_reg[40]_i_1_n_9 ,\frame_64_good_reg[40]_i_1_n_10 ,\frame_64_good_reg[40]_i_1_n_11 ,\frame_64_good_reg[40]_i_1_n_12 ,\frame_64_good_reg[40]_i_1_n_13 ,\frame_64_good_reg[40]_i_1_n_14 ,\frame_64_good_reg[40]_i_1_n_15 }),
        .S(frame_64_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_14 ),
        .Q(frame_64_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_13 ),
        .Q(frame_64_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_12 ),
        .Q(frame_64_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_11 ),
        .Q(frame_64_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_10 ),
        .Q(frame_64_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_9 ),
        .Q(frame_64_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[40]_i_1_n_8 ),
        .Q(frame_64_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_15 ),
        .Q(frame_64_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[48]_i_1 
       (.CI(\frame_64_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[48]_i_1_n_0 ,\frame_64_good_reg[48]_i_1_n_1 ,\frame_64_good_reg[48]_i_1_n_2 ,\frame_64_good_reg[48]_i_1_n_3 ,\frame_64_good_reg[48]_i_1_n_4 ,\frame_64_good_reg[48]_i_1_n_5 ,\frame_64_good_reg[48]_i_1_n_6 ,\frame_64_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[48]_i_1_n_8 ,\frame_64_good_reg[48]_i_1_n_9 ,\frame_64_good_reg[48]_i_1_n_10 ,\frame_64_good_reg[48]_i_1_n_11 ,\frame_64_good_reg[48]_i_1_n_12 ,\frame_64_good_reg[48]_i_1_n_13 ,\frame_64_good_reg[48]_i_1_n_14 ,\frame_64_good_reg[48]_i_1_n_15 }),
        .S(frame_64_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_14 ),
        .Q(frame_64_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_11 ),
        .Q(frame_64_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_13 ),
        .Q(frame_64_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_12 ),
        .Q(frame_64_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_11 ),
        .Q(frame_64_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_10 ),
        .Q(frame_64_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_9 ),
        .Q(frame_64_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[48]_i_1_n_8 ),
        .Q(frame_64_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_15 ),
        .Q(frame_64_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[56]_i_1 
       (.CI(\frame_64_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_64_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_64_good_reg[56]_i_1_n_1 ,\frame_64_good_reg[56]_i_1_n_2 ,\frame_64_good_reg[56]_i_1_n_3 ,\frame_64_good_reg[56]_i_1_n_4 ,\frame_64_good_reg[56]_i_1_n_5 ,\frame_64_good_reg[56]_i_1_n_6 ,\frame_64_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[56]_i_1_n_8 ,\frame_64_good_reg[56]_i_1_n_9 ,\frame_64_good_reg[56]_i_1_n_10 ,\frame_64_good_reg[56]_i_1_n_11 ,\frame_64_good_reg[56]_i_1_n_12 ,\frame_64_good_reg[56]_i_1_n_13 ,\frame_64_good_reg[56]_i_1_n_14 ,\frame_64_good_reg[56]_i_1_n_15 }),
        .S(frame_64_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_14 ),
        .Q(frame_64_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_13 ),
        .Q(frame_64_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_12 ),
        .Q(frame_64_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_10 ),
        .Q(frame_64_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_11 ),
        .Q(frame_64_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_10 ),
        .Q(frame_64_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_9 ),
        .Q(frame_64_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[56]_i_1_n_8 ),
        .Q(frame_64_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_9 ),
        .Q(frame_64_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[0]_i_1_n_8 ),
        .Q(frame_64_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_15 ),
        .Q(frame_64_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_good_reg[8]_i_1 
       (.CI(\frame_64_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_good_reg[8]_i_1_n_0 ,\frame_64_good_reg[8]_i_1_n_1 ,\frame_64_good_reg[8]_i_1_n_2 ,\frame_64_good_reg[8]_i_1_n_3 ,\frame_64_good_reg[8]_i_1_n_4 ,\frame_64_good_reg[8]_i_1_n_5 ,\frame_64_good_reg[8]_i_1_n_6 ,\frame_64_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_good_reg[8]_i_1_n_8 ,\frame_64_good_reg[8]_i_1_n_9 ,\frame_64_good_reg[8]_i_1_n_10 ,\frame_64_good_reg[8]_i_1_n_11 ,\frame_64_good_reg[8]_i_1_n_12 ,\frame_64_good_reg[8]_i_1_n_13 ,\frame_64_good_reg[8]_i_1_n_14 ,\frame_64_good_reg[8]_i_1_n_15 }),
        .S(frame_64_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[4]),
        .CLR(rst_i),
        .D(\frame_64_good_reg[8]_i_1_n_14 ),
        .Q(frame_64_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_64_transed[0]_i_2 
       (.I0(frame_64_transed_reg[0]),
        .O(\frame_64_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_15 ),
        .Q(frame_64_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[0]_i_1_n_0 ,\frame_64_transed_reg[0]_i_1_n_1 ,\frame_64_transed_reg[0]_i_1_n_2 ,\frame_64_transed_reg[0]_i_1_n_3 ,\frame_64_transed_reg[0]_i_1_n_4 ,\frame_64_transed_reg[0]_i_1_n_5 ,\frame_64_transed_reg[0]_i_1_n_6 ,\frame_64_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_64_transed_reg[0]_i_1_n_8 ,\frame_64_transed_reg[0]_i_1_n_9 ,\frame_64_transed_reg[0]_i_1_n_10 ,\frame_64_transed_reg[0]_i_1_n_11 ,\frame_64_transed_reg[0]_i_1_n_12 ,\frame_64_transed_reg[0]_i_1_n_13 ,\frame_64_transed_reg[0]_i_1_n_14 ,\frame_64_transed_reg[0]_i_1_n_15 }),
        .S({frame_64_transed_reg[7:1],\frame_64_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_13 ),
        .Q(frame_64_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_12 ),
        .Q(frame_64_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_11 ),
        .Q(frame_64_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_10 ),
        .Q(frame_64_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_9 ),
        .Q(frame_64_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_8 ),
        .Q(frame_64_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_15 ),
        .Q(frame_64_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[16]_i_1 
       (.CI(\frame_64_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[16]_i_1_n_0 ,\frame_64_transed_reg[16]_i_1_n_1 ,\frame_64_transed_reg[16]_i_1_n_2 ,\frame_64_transed_reg[16]_i_1_n_3 ,\frame_64_transed_reg[16]_i_1_n_4 ,\frame_64_transed_reg[16]_i_1_n_5 ,\frame_64_transed_reg[16]_i_1_n_6 ,\frame_64_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[16]_i_1_n_8 ,\frame_64_transed_reg[16]_i_1_n_9 ,\frame_64_transed_reg[16]_i_1_n_10 ,\frame_64_transed_reg[16]_i_1_n_11 ,\frame_64_transed_reg[16]_i_1_n_12 ,\frame_64_transed_reg[16]_i_1_n_13 ,\frame_64_transed_reg[16]_i_1_n_14 ,\frame_64_transed_reg[16]_i_1_n_15 }),
        .S(frame_64_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_14 ),
        .Q(frame_64_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_13 ),
        .Q(frame_64_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_12 ),
        .Q(frame_64_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_14 ),
        .Q(frame_64_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_11 ),
        .Q(frame_64_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_10 ),
        .Q(frame_64_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_9 ),
        .Q(frame_64_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[16]_i_1_n_8 ),
        .Q(frame_64_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_15 ),
        .Q(frame_64_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[24]_i_1 
       (.CI(\frame_64_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[24]_i_1_n_0 ,\frame_64_transed_reg[24]_i_1_n_1 ,\frame_64_transed_reg[24]_i_1_n_2 ,\frame_64_transed_reg[24]_i_1_n_3 ,\frame_64_transed_reg[24]_i_1_n_4 ,\frame_64_transed_reg[24]_i_1_n_5 ,\frame_64_transed_reg[24]_i_1_n_6 ,\frame_64_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[24]_i_1_n_8 ,\frame_64_transed_reg[24]_i_1_n_9 ,\frame_64_transed_reg[24]_i_1_n_10 ,\frame_64_transed_reg[24]_i_1_n_11 ,\frame_64_transed_reg[24]_i_1_n_12 ,\frame_64_transed_reg[24]_i_1_n_13 ,\frame_64_transed_reg[24]_i_1_n_14 ,\frame_64_transed_reg[24]_i_1_n_15 }),
        .S(frame_64_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_14 ),
        .Q(frame_64_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_13 ),
        .Q(frame_64_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_12 ),
        .Q(frame_64_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_11 ),
        .Q(frame_64_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_10 ),
        .Q(frame_64_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_13 ),
        .Q(frame_64_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_9 ),
        .Q(frame_64_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[24]_i_1_n_8 ),
        .Q(frame_64_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_15 ),
        .Q(frame_64_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[32]_i_1 
       (.CI(\frame_64_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[32]_i_1_n_0 ,\frame_64_transed_reg[32]_i_1_n_1 ,\frame_64_transed_reg[32]_i_1_n_2 ,\frame_64_transed_reg[32]_i_1_n_3 ,\frame_64_transed_reg[32]_i_1_n_4 ,\frame_64_transed_reg[32]_i_1_n_5 ,\frame_64_transed_reg[32]_i_1_n_6 ,\frame_64_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[32]_i_1_n_8 ,\frame_64_transed_reg[32]_i_1_n_9 ,\frame_64_transed_reg[32]_i_1_n_10 ,\frame_64_transed_reg[32]_i_1_n_11 ,\frame_64_transed_reg[32]_i_1_n_12 ,\frame_64_transed_reg[32]_i_1_n_13 ,\frame_64_transed_reg[32]_i_1_n_14 ,\frame_64_transed_reg[32]_i_1_n_15 }),
        .S(frame_64_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_14 ),
        .Q(frame_64_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_13 ),
        .Q(frame_64_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_12 ),
        .Q(frame_64_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_11 ),
        .Q(frame_64_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_10 ),
        .Q(frame_64_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_9 ),
        .Q(frame_64_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[32]_i_1_n_8 ),
        .Q(frame_64_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_12 ),
        .Q(frame_64_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_15 ),
        .Q(frame_64_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[40]_i_1 
       (.CI(\frame_64_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[40]_i_1_n_0 ,\frame_64_transed_reg[40]_i_1_n_1 ,\frame_64_transed_reg[40]_i_1_n_2 ,\frame_64_transed_reg[40]_i_1_n_3 ,\frame_64_transed_reg[40]_i_1_n_4 ,\frame_64_transed_reg[40]_i_1_n_5 ,\frame_64_transed_reg[40]_i_1_n_6 ,\frame_64_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[40]_i_1_n_8 ,\frame_64_transed_reg[40]_i_1_n_9 ,\frame_64_transed_reg[40]_i_1_n_10 ,\frame_64_transed_reg[40]_i_1_n_11 ,\frame_64_transed_reg[40]_i_1_n_12 ,\frame_64_transed_reg[40]_i_1_n_13 ,\frame_64_transed_reg[40]_i_1_n_14 ,\frame_64_transed_reg[40]_i_1_n_15 }),
        .S(frame_64_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_14 ),
        .Q(frame_64_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_13 ),
        .Q(frame_64_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_12 ),
        .Q(frame_64_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_11 ),
        .Q(frame_64_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_10 ),
        .Q(frame_64_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_9 ),
        .Q(frame_64_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[40]_i_1_n_8 ),
        .Q(frame_64_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_15 ),
        .Q(frame_64_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[48]_i_1 
       (.CI(\frame_64_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[48]_i_1_n_0 ,\frame_64_transed_reg[48]_i_1_n_1 ,\frame_64_transed_reg[48]_i_1_n_2 ,\frame_64_transed_reg[48]_i_1_n_3 ,\frame_64_transed_reg[48]_i_1_n_4 ,\frame_64_transed_reg[48]_i_1_n_5 ,\frame_64_transed_reg[48]_i_1_n_6 ,\frame_64_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[48]_i_1_n_8 ,\frame_64_transed_reg[48]_i_1_n_9 ,\frame_64_transed_reg[48]_i_1_n_10 ,\frame_64_transed_reg[48]_i_1_n_11 ,\frame_64_transed_reg[48]_i_1_n_12 ,\frame_64_transed_reg[48]_i_1_n_13 ,\frame_64_transed_reg[48]_i_1_n_14 ,\frame_64_transed_reg[48]_i_1_n_15 }),
        .S(frame_64_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_14 ),
        .Q(frame_64_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_11 ),
        .Q(frame_64_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_13 ),
        .Q(frame_64_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_12 ),
        .Q(frame_64_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_11 ),
        .Q(frame_64_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_10 ),
        .Q(frame_64_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_9 ),
        .Q(frame_64_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[48]_i_1_n_8 ),
        .Q(frame_64_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_15 ),
        .Q(frame_64_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[56]_i_1 
       (.CI(\frame_64_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_64_transed_reg[56]_i_1_CO_UNCONNECTED [7],\frame_64_transed_reg[56]_i_1_n_1 ,\frame_64_transed_reg[56]_i_1_n_2 ,\frame_64_transed_reg[56]_i_1_n_3 ,\frame_64_transed_reg[56]_i_1_n_4 ,\frame_64_transed_reg[56]_i_1_n_5 ,\frame_64_transed_reg[56]_i_1_n_6 ,\frame_64_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[56]_i_1_n_8 ,\frame_64_transed_reg[56]_i_1_n_9 ,\frame_64_transed_reg[56]_i_1_n_10 ,\frame_64_transed_reg[56]_i_1_n_11 ,\frame_64_transed_reg[56]_i_1_n_12 ,\frame_64_transed_reg[56]_i_1_n_13 ,\frame_64_transed_reg[56]_i_1_n_14 ,\frame_64_transed_reg[56]_i_1_n_15 }),
        .S(frame_64_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_14 ),
        .Q(frame_64_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_13 ),
        .Q(frame_64_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_12 ),
        .Q(frame_64_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_10 ),
        .Q(frame_64_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_11 ),
        .Q(frame_64_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_10 ),
        .Q(frame_64_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_9 ),
        .Q(frame_64_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[56]_i_1_n_8 ),
        .Q(frame_64_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_9 ),
        .Q(frame_64_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[0]_i_1_n_8 ),
        .Q(frame_64_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_15 ),
        .Q(frame_64_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_64_transed_reg[8]_i_1 
       (.CI(\frame_64_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_64_transed_reg[8]_i_1_n_0 ,\frame_64_transed_reg[8]_i_1_n_1 ,\frame_64_transed_reg[8]_i_1_n_2 ,\frame_64_transed_reg[8]_i_1_n_3 ,\frame_64_transed_reg[8]_i_1_n_4 ,\frame_64_transed_reg[8]_i_1_n_5 ,\frame_64_transed_reg[8]_i_1_n_6 ,\frame_64_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_64_transed_reg[8]_i_1_n_8 ,\frame_64_transed_reg[8]_i_1_n_9 ,\frame_64_transed_reg[8]_i_1_n_10 ,\frame_64_transed_reg[8]_i_1_n_11 ,\frame_64_transed_reg[8]_i_1_n_12 ,\frame_64_transed_reg[8]_i_1_n_13 ,\frame_64_transed_reg[8]_i_1_n_14 ,\frame_64_transed_reg[8]_i_1_n_15 }),
        .S(frame_64_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_64_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[6]),
        .CLR(rst_i),
        .D(\frame_64_transed_reg[8]_i_1_n_14 ),
        .Q(frame_64_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_65_127_good[0]_i_2 
       (.I0(frame_65_127_good_reg[0]),
        .O(\frame_65_127_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[0]_i_1_n_0 ,\frame_65_127_good_reg[0]_i_1_n_1 ,\frame_65_127_good_reg[0]_i_1_n_2 ,\frame_65_127_good_reg[0]_i_1_n_3 ,\frame_65_127_good_reg[0]_i_1_n_4 ,\frame_65_127_good_reg[0]_i_1_n_5 ,\frame_65_127_good_reg[0]_i_1_n_6 ,\frame_65_127_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_65_127_good_reg[0]_i_1_n_8 ,\frame_65_127_good_reg[0]_i_1_n_9 ,\frame_65_127_good_reg[0]_i_1_n_10 ,\frame_65_127_good_reg[0]_i_1_n_11 ,\frame_65_127_good_reg[0]_i_1_n_12 ,\frame_65_127_good_reg[0]_i_1_n_13 ,\frame_65_127_good_reg[0]_i_1_n_14 ,\frame_65_127_good_reg[0]_i_1_n_15 }),
        .S({frame_65_127_good_reg[7:1],\frame_65_127_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[16]_i_1 
       (.CI(\frame_65_127_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[16]_i_1_n_0 ,\frame_65_127_good_reg[16]_i_1_n_1 ,\frame_65_127_good_reg[16]_i_1_n_2 ,\frame_65_127_good_reg[16]_i_1_n_3 ,\frame_65_127_good_reg[16]_i_1_n_4 ,\frame_65_127_good_reg[16]_i_1_n_5 ,\frame_65_127_good_reg[16]_i_1_n_6 ,\frame_65_127_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[16]_i_1_n_8 ,\frame_65_127_good_reg[16]_i_1_n_9 ,\frame_65_127_good_reg[16]_i_1_n_10 ,\frame_65_127_good_reg[16]_i_1_n_11 ,\frame_65_127_good_reg[16]_i_1_n_12 ,\frame_65_127_good_reg[16]_i_1_n_13 ,\frame_65_127_good_reg[16]_i_1_n_14 ,\frame_65_127_good_reg[16]_i_1_n_15 }),
        .S(frame_65_127_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[16]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[24]_i_1 
       (.CI(\frame_65_127_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[24]_i_1_n_0 ,\frame_65_127_good_reg[24]_i_1_n_1 ,\frame_65_127_good_reg[24]_i_1_n_2 ,\frame_65_127_good_reg[24]_i_1_n_3 ,\frame_65_127_good_reg[24]_i_1_n_4 ,\frame_65_127_good_reg[24]_i_1_n_5 ,\frame_65_127_good_reg[24]_i_1_n_6 ,\frame_65_127_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[24]_i_1_n_8 ,\frame_65_127_good_reg[24]_i_1_n_9 ,\frame_65_127_good_reg[24]_i_1_n_10 ,\frame_65_127_good_reg[24]_i_1_n_11 ,\frame_65_127_good_reg[24]_i_1_n_12 ,\frame_65_127_good_reg[24]_i_1_n_13 ,\frame_65_127_good_reg[24]_i_1_n_14 ,\frame_65_127_good_reg[24]_i_1_n_15 }),
        .S(frame_65_127_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[24]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[32]_i_1 
       (.CI(\frame_65_127_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[32]_i_1_n_0 ,\frame_65_127_good_reg[32]_i_1_n_1 ,\frame_65_127_good_reg[32]_i_1_n_2 ,\frame_65_127_good_reg[32]_i_1_n_3 ,\frame_65_127_good_reg[32]_i_1_n_4 ,\frame_65_127_good_reg[32]_i_1_n_5 ,\frame_65_127_good_reg[32]_i_1_n_6 ,\frame_65_127_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[32]_i_1_n_8 ,\frame_65_127_good_reg[32]_i_1_n_9 ,\frame_65_127_good_reg[32]_i_1_n_10 ,\frame_65_127_good_reg[32]_i_1_n_11 ,\frame_65_127_good_reg[32]_i_1_n_12 ,\frame_65_127_good_reg[32]_i_1_n_13 ,\frame_65_127_good_reg[32]_i_1_n_14 ,\frame_65_127_good_reg[32]_i_1_n_15 }),
        .S(frame_65_127_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[32]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[40]_i_1 
       (.CI(\frame_65_127_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[40]_i_1_n_0 ,\frame_65_127_good_reg[40]_i_1_n_1 ,\frame_65_127_good_reg[40]_i_1_n_2 ,\frame_65_127_good_reg[40]_i_1_n_3 ,\frame_65_127_good_reg[40]_i_1_n_4 ,\frame_65_127_good_reg[40]_i_1_n_5 ,\frame_65_127_good_reg[40]_i_1_n_6 ,\frame_65_127_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[40]_i_1_n_8 ,\frame_65_127_good_reg[40]_i_1_n_9 ,\frame_65_127_good_reg[40]_i_1_n_10 ,\frame_65_127_good_reg[40]_i_1_n_11 ,\frame_65_127_good_reg[40]_i_1_n_12 ,\frame_65_127_good_reg[40]_i_1_n_13 ,\frame_65_127_good_reg[40]_i_1_n_14 ,\frame_65_127_good_reg[40]_i_1_n_15 }),
        .S(frame_65_127_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[40]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[48]_i_1 
       (.CI(\frame_65_127_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[48]_i_1_n_0 ,\frame_65_127_good_reg[48]_i_1_n_1 ,\frame_65_127_good_reg[48]_i_1_n_2 ,\frame_65_127_good_reg[48]_i_1_n_3 ,\frame_65_127_good_reg[48]_i_1_n_4 ,\frame_65_127_good_reg[48]_i_1_n_5 ,\frame_65_127_good_reg[48]_i_1_n_6 ,\frame_65_127_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[48]_i_1_n_8 ,\frame_65_127_good_reg[48]_i_1_n_9 ,\frame_65_127_good_reg[48]_i_1_n_10 ,\frame_65_127_good_reg[48]_i_1_n_11 ,\frame_65_127_good_reg[48]_i_1_n_12 ,\frame_65_127_good_reg[48]_i_1_n_13 ,\frame_65_127_good_reg[48]_i_1_n_14 ,\frame_65_127_good_reg[48]_i_1_n_15 }),
        .S(frame_65_127_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[48]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[56]_i_1 
       (.CI(\frame_65_127_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_65_127_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_65_127_good_reg[56]_i_1_n_1 ,\frame_65_127_good_reg[56]_i_1_n_2 ,\frame_65_127_good_reg[56]_i_1_n_3 ,\frame_65_127_good_reg[56]_i_1_n_4 ,\frame_65_127_good_reg[56]_i_1_n_5 ,\frame_65_127_good_reg[56]_i_1_n_6 ,\frame_65_127_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[56]_i_1_n_8 ,\frame_65_127_good_reg[56]_i_1_n_9 ,\frame_65_127_good_reg[56]_i_1_n_10 ,\frame_65_127_good_reg[56]_i_1_n_11 ,\frame_65_127_good_reg[56]_i_1_n_12 ,\frame_65_127_good_reg[56]_i_1_n_13 ,\frame_65_127_good_reg[56]_i_1_n_14 ,\frame_65_127_good_reg[56]_i_1_n_15 }),
        .S(frame_65_127_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_13 ),
        .Q(frame_65_127_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_12 ),
        .Q(frame_65_127_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_11 ),
        .Q(frame_65_127_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_10 ),
        .Q(frame_65_127_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[56]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_9 ),
        .Q(frame_65_127_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[0]_i_1_n_8 ),
        .Q(frame_65_127_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_15 ),
        .Q(frame_65_127_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_good_reg[8]_i_1 
       (.CI(\frame_65_127_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_good_reg[8]_i_1_n_0 ,\frame_65_127_good_reg[8]_i_1_n_1 ,\frame_65_127_good_reg[8]_i_1_n_2 ,\frame_65_127_good_reg[8]_i_1_n_3 ,\frame_65_127_good_reg[8]_i_1_n_4 ,\frame_65_127_good_reg[8]_i_1_n_5 ,\frame_65_127_good_reg[8]_i_1_n_6 ,\frame_65_127_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_good_reg[8]_i_1_n_8 ,\frame_65_127_good_reg[8]_i_1_n_9 ,\frame_65_127_good_reg[8]_i_1_n_10 ,\frame_65_127_good_reg[8]_i_1_n_11 ,\frame_65_127_good_reg[8]_i_1_n_12 ,\frame_65_127_good_reg[8]_i_1_n_13 ,\frame_65_127_good_reg[8]_i_1_n_14 ,\frame_65_127_good_reg[8]_i_1_n_15 }),
        .S(frame_65_127_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[5]),
        .CLR(rst_i),
        .D(\frame_65_127_good_reg[8]_i_1_n_14 ),
        .Q(frame_65_127_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_65_127_transed[0]_i_2 
       (.I0(frame_65_127_transed_reg[0]),
        .O(\frame_65_127_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[0]_i_1_n_0 ,\frame_65_127_transed_reg[0]_i_1_n_1 ,\frame_65_127_transed_reg[0]_i_1_n_2 ,\frame_65_127_transed_reg[0]_i_1_n_3 ,\frame_65_127_transed_reg[0]_i_1_n_4 ,\frame_65_127_transed_reg[0]_i_1_n_5 ,\frame_65_127_transed_reg[0]_i_1_n_6 ,\frame_65_127_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_65_127_transed_reg[0]_i_1_n_8 ,\frame_65_127_transed_reg[0]_i_1_n_9 ,\frame_65_127_transed_reg[0]_i_1_n_10 ,\frame_65_127_transed_reg[0]_i_1_n_11 ,\frame_65_127_transed_reg[0]_i_1_n_12 ,\frame_65_127_transed_reg[0]_i_1_n_13 ,\frame_65_127_transed_reg[0]_i_1_n_14 ,\frame_65_127_transed_reg[0]_i_1_n_15 }),
        .S({frame_65_127_transed_reg[7:1],\frame_65_127_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[16]_i_1 
       (.CI(\frame_65_127_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[16]_i_1_n_0 ,\frame_65_127_transed_reg[16]_i_1_n_1 ,\frame_65_127_transed_reg[16]_i_1_n_2 ,\frame_65_127_transed_reg[16]_i_1_n_3 ,\frame_65_127_transed_reg[16]_i_1_n_4 ,\frame_65_127_transed_reg[16]_i_1_n_5 ,\frame_65_127_transed_reg[16]_i_1_n_6 ,\frame_65_127_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[16]_i_1_n_8 ,\frame_65_127_transed_reg[16]_i_1_n_9 ,\frame_65_127_transed_reg[16]_i_1_n_10 ,\frame_65_127_transed_reg[16]_i_1_n_11 ,\frame_65_127_transed_reg[16]_i_1_n_12 ,\frame_65_127_transed_reg[16]_i_1_n_13 ,\frame_65_127_transed_reg[16]_i_1_n_14 ,\frame_65_127_transed_reg[16]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[16]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[24]_i_1 
       (.CI(\frame_65_127_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[24]_i_1_n_0 ,\frame_65_127_transed_reg[24]_i_1_n_1 ,\frame_65_127_transed_reg[24]_i_1_n_2 ,\frame_65_127_transed_reg[24]_i_1_n_3 ,\frame_65_127_transed_reg[24]_i_1_n_4 ,\frame_65_127_transed_reg[24]_i_1_n_5 ,\frame_65_127_transed_reg[24]_i_1_n_6 ,\frame_65_127_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[24]_i_1_n_8 ,\frame_65_127_transed_reg[24]_i_1_n_9 ,\frame_65_127_transed_reg[24]_i_1_n_10 ,\frame_65_127_transed_reg[24]_i_1_n_11 ,\frame_65_127_transed_reg[24]_i_1_n_12 ,\frame_65_127_transed_reg[24]_i_1_n_13 ,\frame_65_127_transed_reg[24]_i_1_n_14 ,\frame_65_127_transed_reg[24]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[24]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[32]_i_1 
       (.CI(\frame_65_127_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[32]_i_1_n_0 ,\frame_65_127_transed_reg[32]_i_1_n_1 ,\frame_65_127_transed_reg[32]_i_1_n_2 ,\frame_65_127_transed_reg[32]_i_1_n_3 ,\frame_65_127_transed_reg[32]_i_1_n_4 ,\frame_65_127_transed_reg[32]_i_1_n_5 ,\frame_65_127_transed_reg[32]_i_1_n_6 ,\frame_65_127_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[32]_i_1_n_8 ,\frame_65_127_transed_reg[32]_i_1_n_9 ,\frame_65_127_transed_reg[32]_i_1_n_10 ,\frame_65_127_transed_reg[32]_i_1_n_11 ,\frame_65_127_transed_reg[32]_i_1_n_12 ,\frame_65_127_transed_reg[32]_i_1_n_13 ,\frame_65_127_transed_reg[32]_i_1_n_14 ,\frame_65_127_transed_reg[32]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[32]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[40]_i_1 
       (.CI(\frame_65_127_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[40]_i_1_n_0 ,\frame_65_127_transed_reg[40]_i_1_n_1 ,\frame_65_127_transed_reg[40]_i_1_n_2 ,\frame_65_127_transed_reg[40]_i_1_n_3 ,\frame_65_127_transed_reg[40]_i_1_n_4 ,\frame_65_127_transed_reg[40]_i_1_n_5 ,\frame_65_127_transed_reg[40]_i_1_n_6 ,\frame_65_127_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[40]_i_1_n_8 ,\frame_65_127_transed_reg[40]_i_1_n_9 ,\frame_65_127_transed_reg[40]_i_1_n_10 ,\frame_65_127_transed_reg[40]_i_1_n_11 ,\frame_65_127_transed_reg[40]_i_1_n_12 ,\frame_65_127_transed_reg[40]_i_1_n_13 ,\frame_65_127_transed_reg[40]_i_1_n_14 ,\frame_65_127_transed_reg[40]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[40]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[48]_i_1 
       (.CI(\frame_65_127_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[48]_i_1_n_0 ,\frame_65_127_transed_reg[48]_i_1_n_1 ,\frame_65_127_transed_reg[48]_i_1_n_2 ,\frame_65_127_transed_reg[48]_i_1_n_3 ,\frame_65_127_transed_reg[48]_i_1_n_4 ,\frame_65_127_transed_reg[48]_i_1_n_5 ,\frame_65_127_transed_reg[48]_i_1_n_6 ,\frame_65_127_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[48]_i_1_n_8 ,\frame_65_127_transed_reg[48]_i_1_n_9 ,\frame_65_127_transed_reg[48]_i_1_n_10 ,\frame_65_127_transed_reg[48]_i_1_n_11 ,\frame_65_127_transed_reg[48]_i_1_n_12 ,\frame_65_127_transed_reg[48]_i_1_n_13 ,\frame_65_127_transed_reg[48]_i_1_n_14 ,\frame_65_127_transed_reg[48]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[48]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[56]_i_1 
       (.CI(\frame_65_127_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_65_127_transed_reg[56]_i_1_CO_UNCONNECTED [7],\frame_65_127_transed_reg[56]_i_1_n_1 ,\frame_65_127_transed_reg[56]_i_1_n_2 ,\frame_65_127_transed_reg[56]_i_1_n_3 ,\frame_65_127_transed_reg[56]_i_1_n_4 ,\frame_65_127_transed_reg[56]_i_1_n_5 ,\frame_65_127_transed_reg[56]_i_1_n_6 ,\frame_65_127_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[56]_i_1_n_8 ,\frame_65_127_transed_reg[56]_i_1_n_9 ,\frame_65_127_transed_reg[56]_i_1_n_10 ,\frame_65_127_transed_reg[56]_i_1_n_11 ,\frame_65_127_transed_reg[56]_i_1_n_12 ,\frame_65_127_transed_reg[56]_i_1_n_13 ,\frame_65_127_transed_reg[56]_i_1_n_14 ,\frame_65_127_transed_reg[56]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_13 ),
        .Q(frame_65_127_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_12 ),
        .Q(frame_65_127_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_11 ),
        .Q(frame_65_127_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_10 ),
        .Q(frame_65_127_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[56]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_9 ),
        .Q(frame_65_127_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[0]_i_1_n_8 ),
        .Q(frame_65_127_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_15 ),
        .Q(frame_65_127_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_65_127_transed_reg[8]_i_1 
       (.CI(\frame_65_127_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_65_127_transed_reg[8]_i_1_n_0 ,\frame_65_127_transed_reg[8]_i_1_n_1 ,\frame_65_127_transed_reg[8]_i_1_n_2 ,\frame_65_127_transed_reg[8]_i_1_n_3 ,\frame_65_127_transed_reg[8]_i_1_n_4 ,\frame_65_127_transed_reg[8]_i_1_n_5 ,\frame_65_127_transed_reg[8]_i_1_n_6 ,\frame_65_127_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_65_127_transed_reg[8]_i_1_n_8 ,\frame_65_127_transed_reg[8]_i_1_n_9 ,\frame_65_127_transed_reg[8]_i_1_n_10 ,\frame_65_127_transed_reg[8]_i_1_n_11 ,\frame_65_127_transed_reg[8]_i_1_n_12 ,\frame_65_127_transed_reg[8]_i_1_n_13 ,\frame_65_127_transed_reg[8]_i_1_n_14 ,\frame_65_127_transed_reg[8]_i_1_n_15 }),
        .S(frame_65_127_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_65_127_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[7]),
        .CLR(rst_i),
        .D(\frame_65_127_transed_reg[8]_i_1_n_14 ),
        .Q(frame_65_127_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \frame_received_good[0]_i_2 
       (.I0(frame_received_good_reg[0]),
        .O(\frame_received_good[0]_i_2_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \frame_received_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .D(\frame_received_good_reg[0]_i_1_n_15 ),
        .PRE(rst_i),
        .Q(frame_received_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[0]_i_1_n_0 ,\frame_received_good_reg[0]_i_1_n_1 ,\frame_received_good_reg[0]_i_1_n_2 ,\frame_received_good_reg[0]_i_1_n_3 ,\frame_received_good_reg[0]_i_1_n_4 ,\frame_received_good_reg[0]_i_1_n_5 ,\frame_received_good_reg[0]_i_1_n_6 ,\frame_received_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\frame_received_good_reg[0]_i_1_n_8 ,\frame_received_good_reg[0]_i_1_n_9 ,\frame_received_good_reg[0]_i_1_n_10 ,\frame_received_good_reg[0]_i_1_n_11 ,\frame_received_good_reg[0]_i_1_n_12 ,\frame_received_good_reg[0]_i_1_n_13 ,\frame_received_good_reg[0]_i_1_n_14 ,\frame_received_good_reg[0]_i_1_n_15 }),
        .S({frame_received_good_reg[7:1],\frame_received_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_13 ),
        .Q(frame_received_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_12 ),
        .Q(frame_received_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_11 ),
        .Q(frame_received_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_10 ),
        .Q(frame_received_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_9 ),
        .Q(frame_received_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_8 ),
        .Q(frame_received_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_15 ),
        .Q(frame_received_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[16]_i_1 
       (.CI(\frame_received_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[16]_i_1_n_0 ,\frame_received_good_reg[16]_i_1_n_1 ,\frame_received_good_reg[16]_i_1_n_2 ,\frame_received_good_reg[16]_i_1_n_3 ,\frame_received_good_reg[16]_i_1_n_4 ,\frame_received_good_reg[16]_i_1_n_5 ,\frame_received_good_reg[16]_i_1_n_6 ,\frame_received_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[16]_i_1_n_8 ,\frame_received_good_reg[16]_i_1_n_9 ,\frame_received_good_reg[16]_i_1_n_10 ,\frame_received_good_reg[16]_i_1_n_11 ,\frame_received_good_reg[16]_i_1_n_12 ,\frame_received_good_reg[16]_i_1_n_13 ,\frame_received_good_reg[16]_i_1_n_14 ,\frame_received_good_reg[16]_i_1_n_15 }),
        .S(frame_received_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_14 ),
        .Q(frame_received_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_13 ),
        .Q(frame_received_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_12 ),
        .Q(frame_received_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_14 ),
        .Q(frame_received_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_11 ),
        .Q(frame_received_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_10 ),
        .Q(frame_received_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_9 ),
        .Q(frame_received_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[16]_i_1_n_8 ),
        .Q(frame_received_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_15 ),
        .Q(frame_received_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[24]_i_1 
       (.CI(\frame_received_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[24]_i_1_n_0 ,\frame_received_good_reg[24]_i_1_n_1 ,\frame_received_good_reg[24]_i_1_n_2 ,\frame_received_good_reg[24]_i_1_n_3 ,\frame_received_good_reg[24]_i_1_n_4 ,\frame_received_good_reg[24]_i_1_n_5 ,\frame_received_good_reg[24]_i_1_n_6 ,\frame_received_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[24]_i_1_n_8 ,\frame_received_good_reg[24]_i_1_n_9 ,\frame_received_good_reg[24]_i_1_n_10 ,\frame_received_good_reg[24]_i_1_n_11 ,\frame_received_good_reg[24]_i_1_n_12 ,\frame_received_good_reg[24]_i_1_n_13 ,\frame_received_good_reg[24]_i_1_n_14 ,\frame_received_good_reg[24]_i_1_n_15 }),
        .S(frame_received_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_14 ),
        .Q(frame_received_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_13 ),
        .Q(frame_received_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_12 ),
        .Q(frame_received_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_11 ),
        .Q(frame_received_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_10 ),
        .Q(frame_received_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_13 ),
        .Q(frame_received_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_9 ),
        .Q(frame_received_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[24]_i_1_n_8 ),
        .Q(frame_received_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_15 ),
        .Q(frame_received_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[32]_i_1 
       (.CI(\frame_received_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[32]_i_1_n_0 ,\frame_received_good_reg[32]_i_1_n_1 ,\frame_received_good_reg[32]_i_1_n_2 ,\frame_received_good_reg[32]_i_1_n_3 ,\frame_received_good_reg[32]_i_1_n_4 ,\frame_received_good_reg[32]_i_1_n_5 ,\frame_received_good_reg[32]_i_1_n_6 ,\frame_received_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[32]_i_1_n_8 ,\frame_received_good_reg[32]_i_1_n_9 ,\frame_received_good_reg[32]_i_1_n_10 ,\frame_received_good_reg[32]_i_1_n_11 ,\frame_received_good_reg[32]_i_1_n_12 ,\frame_received_good_reg[32]_i_1_n_13 ,\frame_received_good_reg[32]_i_1_n_14 ,\frame_received_good_reg[32]_i_1_n_15 }),
        .S(frame_received_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_14 ),
        .Q(frame_received_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_13 ),
        .Q(frame_received_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_12 ),
        .Q(frame_received_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_11 ),
        .Q(frame_received_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_10 ),
        .Q(frame_received_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_9 ),
        .Q(frame_received_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[32]_i_1_n_8 ),
        .Q(frame_received_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_12 ),
        .Q(frame_received_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_15 ),
        .Q(frame_received_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[40]_i_1 
       (.CI(\frame_received_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[40]_i_1_n_0 ,\frame_received_good_reg[40]_i_1_n_1 ,\frame_received_good_reg[40]_i_1_n_2 ,\frame_received_good_reg[40]_i_1_n_3 ,\frame_received_good_reg[40]_i_1_n_4 ,\frame_received_good_reg[40]_i_1_n_5 ,\frame_received_good_reg[40]_i_1_n_6 ,\frame_received_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[40]_i_1_n_8 ,\frame_received_good_reg[40]_i_1_n_9 ,\frame_received_good_reg[40]_i_1_n_10 ,\frame_received_good_reg[40]_i_1_n_11 ,\frame_received_good_reg[40]_i_1_n_12 ,\frame_received_good_reg[40]_i_1_n_13 ,\frame_received_good_reg[40]_i_1_n_14 ,\frame_received_good_reg[40]_i_1_n_15 }),
        .S(frame_received_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_14 ),
        .Q(frame_received_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_13 ),
        .Q(frame_received_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_12 ),
        .Q(frame_received_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_11 ),
        .Q(frame_received_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_10 ),
        .Q(frame_received_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_9 ),
        .Q(frame_received_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[40]_i_1_n_8 ),
        .Q(frame_received_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_15 ),
        .Q(frame_received_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[48]_i_1 
       (.CI(\frame_received_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[48]_i_1_n_0 ,\frame_received_good_reg[48]_i_1_n_1 ,\frame_received_good_reg[48]_i_1_n_2 ,\frame_received_good_reg[48]_i_1_n_3 ,\frame_received_good_reg[48]_i_1_n_4 ,\frame_received_good_reg[48]_i_1_n_5 ,\frame_received_good_reg[48]_i_1_n_6 ,\frame_received_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[48]_i_1_n_8 ,\frame_received_good_reg[48]_i_1_n_9 ,\frame_received_good_reg[48]_i_1_n_10 ,\frame_received_good_reg[48]_i_1_n_11 ,\frame_received_good_reg[48]_i_1_n_12 ,\frame_received_good_reg[48]_i_1_n_13 ,\frame_received_good_reg[48]_i_1_n_14 ,\frame_received_good_reg[48]_i_1_n_15 }),
        .S(frame_received_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_14 ),
        .Q(frame_received_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_11 ),
        .Q(frame_received_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_13 ),
        .Q(frame_received_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_12 ),
        .Q(frame_received_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_11 ),
        .Q(frame_received_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_10 ),
        .Q(frame_received_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_9 ),
        .Q(frame_received_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[48]_i_1_n_8 ),
        .Q(frame_received_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_15 ),
        .Q(frame_received_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[56]_i_1 
       (.CI(\frame_received_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_frame_received_good_reg[56]_i_1_CO_UNCONNECTED [7],\frame_received_good_reg[56]_i_1_n_1 ,\frame_received_good_reg[56]_i_1_n_2 ,\frame_received_good_reg[56]_i_1_n_3 ,\frame_received_good_reg[56]_i_1_n_4 ,\frame_received_good_reg[56]_i_1_n_5 ,\frame_received_good_reg[56]_i_1_n_6 ,\frame_received_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[56]_i_1_n_8 ,\frame_received_good_reg[56]_i_1_n_9 ,\frame_received_good_reg[56]_i_1_n_10 ,\frame_received_good_reg[56]_i_1_n_11 ,\frame_received_good_reg[56]_i_1_n_12 ,\frame_received_good_reg[56]_i_1_n_13 ,\frame_received_good_reg[56]_i_1_n_14 ,\frame_received_good_reg[56]_i_1_n_15 }),
        .S(frame_received_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_14 ),
        .Q(frame_received_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_13 ),
        .Q(frame_received_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_12 ),
        .Q(frame_received_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_10 ),
        .Q(frame_received_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_11 ),
        .Q(frame_received_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_10 ),
        .Q(frame_received_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_9 ),
        .Q(frame_received_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[56]_i_1_n_8 ),
        .Q(frame_received_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_9 ),
        .Q(frame_received_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[0]_i_1_n_8 ),
        .Q(frame_received_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_15 ),
        .Q(frame_received_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \frame_received_good_reg[8]_i_1 
       (.CI(\frame_received_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\frame_received_good_reg[8]_i_1_n_0 ,\frame_received_good_reg[8]_i_1_n_1 ,\frame_received_good_reg[8]_i_1_n_2 ,\frame_received_good_reg[8]_i_1_n_3 ,\frame_received_good_reg[8]_i_1_n_4 ,\frame_received_good_reg[8]_i_1_n_5 ,\frame_received_good_reg[8]_i_1_n_6 ,\frame_received_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\frame_received_good_reg[8]_i_1_n_8 ,\frame_received_good_reg[8]_i_1_n_9 ,\frame_received_good_reg[8]_i_1_n_10 ,\frame_received_good_reg[8]_i_1_n_11 ,\frame_received_good_reg[8]_i_1_n_12 ,\frame_received_good_reg[8]_i_1_n_13 ,\frame_received_good_reg[8]_i_1_n_14 ,\frame_received_good_reg[8]_i_1_n_15 }),
        .S(frame_received_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \frame_received_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[0]),
        .CLR(rst_i),
        .D(\frame_received_good_reg[8]_i_1_n_14 ),
        .Q(frame_received_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \good_frame_transed[0]_i_2 
       (.I0(good_frame_transed_reg[0]),
        .O(\good_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_15 ),
        .Q(good_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[0]_i_1_n_0 ,\good_frame_transed_reg[0]_i_1_n_1 ,\good_frame_transed_reg[0]_i_1_n_2 ,\good_frame_transed_reg[0]_i_1_n_3 ,\good_frame_transed_reg[0]_i_1_n_4 ,\good_frame_transed_reg[0]_i_1_n_5 ,\good_frame_transed_reg[0]_i_1_n_6 ,\good_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\good_frame_transed_reg[0]_i_1_n_8 ,\good_frame_transed_reg[0]_i_1_n_9 ,\good_frame_transed_reg[0]_i_1_n_10 ,\good_frame_transed_reg[0]_i_1_n_11 ,\good_frame_transed_reg[0]_i_1_n_12 ,\good_frame_transed_reg[0]_i_1_n_13 ,\good_frame_transed_reg[0]_i_1_n_14 ,\good_frame_transed_reg[0]_i_1_n_15 }),
        .S({good_frame_transed_reg[7:1],\good_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_13 ),
        .Q(good_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_12 ),
        .Q(good_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_11 ),
        .Q(good_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_10 ),
        .Q(good_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_9 ),
        .Q(good_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_8 ),
        .Q(good_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_15 ),
        .Q(good_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[16]_i_1 
       (.CI(\good_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[16]_i_1_n_0 ,\good_frame_transed_reg[16]_i_1_n_1 ,\good_frame_transed_reg[16]_i_1_n_2 ,\good_frame_transed_reg[16]_i_1_n_3 ,\good_frame_transed_reg[16]_i_1_n_4 ,\good_frame_transed_reg[16]_i_1_n_5 ,\good_frame_transed_reg[16]_i_1_n_6 ,\good_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[16]_i_1_n_8 ,\good_frame_transed_reg[16]_i_1_n_9 ,\good_frame_transed_reg[16]_i_1_n_10 ,\good_frame_transed_reg[16]_i_1_n_11 ,\good_frame_transed_reg[16]_i_1_n_12 ,\good_frame_transed_reg[16]_i_1_n_13 ,\good_frame_transed_reg[16]_i_1_n_14 ,\good_frame_transed_reg[16]_i_1_n_15 }),
        .S(good_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_14 ),
        .Q(good_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_13 ),
        .Q(good_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_12 ),
        .Q(good_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_14 ),
        .Q(good_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_11 ),
        .Q(good_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_10 ),
        .Q(good_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_9 ),
        .Q(good_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[16]_i_1_n_8 ),
        .Q(good_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_15 ),
        .Q(good_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[24]_i_1 
       (.CI(\good_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[24]_i_1_n_0 ,\good_frame_transed_reg[24]_i_1_n_1 ,\good_frame_transed_reg[24]_i_1_n_2 ,\good_frame_transed_reg[24]_i_1_n_3 ,\good_frame_transed_reg[24]_i_1_n_4 ,\good_frame_transed_reg[24]_i_1_n_5 ,\good_frame_transed_reg[24]_i_1_n_6 ,\good_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[24]_i_1_n_8 ,\good_frame_transed_reg[24]_i_1_n_9 ,\good_frame_transed_reg[24]_i_1_n_10 ,\good_frame_transed_reg[24]_i_1_n_11 ,\good_frame_transed_reg[24]_i_1_n_12 ,\good_frame_transed_reg[24]_i_1_n_13 ,\good_frame_transed_reg[24]_i_1_n_14 ,\good_frame_transed_reg[24]_i_1_n_15 }),
        .S(good_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_14 ),
        .Q(good_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_13 ),
        .Q(good_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_12 ),
        .Q(good_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_11 ),
        .Q(good_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_10 ),
        .Q(good_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_13 ),
        .Q(good_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_9 ),
        .Q(good_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[24]_i_1_n_8 ),
        .Q(good_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_15 ),
        .Q(good_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[32]_i_1 
       (.CI(\good_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[32]_i_1_n_0 ,\good_frame_transed_reg[32]_i_1_n_1 ,\good_frame_transed_reg[32]_i_1_n_2 ,\good_frame_transed_reg[32]_i_1_n_3 ,\good_frame_transed_reg[32]_i_1_n_4 ,\good_frame_transed_reg[32]_i_1_n_5 ,\good_frame_transed_reg[32]_i_1_n_6 ,\good_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[32]_i_1_n_8 ,\good_frame_transed_reg[32]_i_1_n_9 ,\good_frame_transed_reg[32]_i_1_n_10 ,\good_frame_transed_reg[32]_i_1_n_11 ,\good_frame_transed_reg[32]_i_1_n_12 ,\good_frame_transed_reg[32]_i_1_n_13 ,\good_frame_transed_reg[32]_i_1_n_14 ,\good_frame_transed_reg[32]_i_1_n_15 }),
        .S(good_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_14 ),
        .Q(good_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_13 ),
        .Q(good_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_12 ),
        .Q(good_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_11 ),
        .Q(good_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_10 ),
        .Q(good_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_9 ),
        .Q(good_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[32]_i_1_n_8 ),
        .Q(good_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_12 ),
        .Q(good_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_15 ),
        .Q(good_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[40]_i_1 
       (.CI(\good_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[40]_i_1_n_0 ,\good_frame_transed_reg[40]_i_1_n_1 ,\good_frame_transed_reg[40]_i_1_n_2 ,\good_frame_transed_reg[40]_i_1_n_3 ,\good_frame_transed_reg[40]_i_1_n_4 ,\good_frame_transed_reg[40]_i_1_n_5 ,\good_frame_transed_reg[40]_i_1_n_6 ,\good_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[40]_i_1_n_8 ,\good_frame_transed_reg[40]_i_1_n_9 ,\good_frame_transed_reg[40]_i_1_n_10 ,\good_frame_transed_reg[40]_i_1_n_11 ,\good_frame_transed_reg[40]_i_1_n_12 ,\good_frame_transed_reg[40]_i_1_n_13 ,\good_frame_transed_reg[40]_i_1_n_14 ,\good_frame_transed_reg[40]_i_1_n_15 }),
        .S(good_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_14 ),
        .Q(good_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_13 ),
        .Q(good_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_12 ),
        .Q(good_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_11 ),
        .Q(good_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_10 ),
        .Q(good_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_9 ),
        .Q(good_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[40]_i_1_n_8 ),
        .Q(good_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_15 ),
        .Q(good_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[48]_i_1 
       (.CI(\good_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[48]_i_1_n_0 ,\good_frame_transed_reg[48]_i_1_n_1 ,\good_frame_transed_reg[48]_i_1_n_2 ,\good_frame_transed_reg[48]_i_1_n_3 ,\good_frame_transed_reg[48]_i_1_n_4 ,\good_frame_transed_reg[48]_i_1_n_5 ,\good_frame_transed_reg[48]_i_1_n_6 ,\good_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[48]_i_1_n_8 ,\good_frame_transed_reg[48]_i_1_n_9 ,\good_frame_transed_reg[48]_i_1_n_10 ,\good_frame_transed_reg[48]_i_1_n_11 ,\good_frame_transed_reg[48]_i_1_n_12 ,\good_frame_transed_reg[48]_i_1_n_13 ,\good_frame_transed_reg[48]_i_1_n_14 ,\good_frame_transed_reg[48]_i_1_n_15 }),
        .S(good_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_14 ),
        .Q(good_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_11 ),
        .Q(good_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_13 ),
        .Q(good_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_12 ),
        .Q(good_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_11 ),
        .Q(good_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_10 ),
        .Q(good_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_9 ),
        .Q(good_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[48]_i_1_n_8 ),
        .Q(good_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_15 ),
        .Q(good_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[56]_i_1 
       (.CI(\good_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_good_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\good_frame_transed_reg[56]_i_1_n_1 ,\good_frame_transed_reg[56]_i_1_n_2 ,\good_frame_transed_reg[56]_i_1_n_3 ,\good_frame_transed_reg[56]_i_1_n_4 ,\good_frame_transed_reg[56]_i_1_n_5 ,\good_frame_transed_reg[56]_i_1_n_6 ,\good_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[56]_i_1_n_8 ,\good_frame_transed_reg[56]_i_1_n_9 ,\good_frame_transed_reg[56]_i_1_n_10 ,\good_frame_transed_reg[56]_i_1_n_11 ,\good_frame_transed_reg[56]_i_1_n_12 ,\good_frame_transed_reg[56]_i_1_n_13 ,\good_frame_transed_reg[56]_i_1_n_14 ,\good_frame_transed_reg[56]_i_1_n_15 }),
        .S(good_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_14 ),
        .Q(good_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_13 ),
        .Q(good_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_12 ),
        .Q(good_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_10 ),
        .Q(good_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_11 ),
        .Q(good_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_10 ),
        .Q(good_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_9 ),
        .Q(good_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[56]_i_1_n_8 ),
        .Q(good_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_9 ),
        .Q(good_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[0]_i_1_n_8 ),
        .Q(good_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_15 ),
        .Q(good_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \good_frame_transed_reg[8]_i_1 
       (.CI(\good_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\good_frame_transed_reg[8]_i_1_n_0 ,\good_frame_transed_reg[8]_i_1_n_1 ,\good_frame_transed_reg[8]_i_1_n_2 ,\good_frame_transed_reg[8]_i_1_n_3 ,\good_frame_transed_reg[8]_i_1_n_4 ,\good_frame_transed_reg[8]_i_1_n_5 ,\good_frame_transed_reg[8]_i_1_n_6 ,\good_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\good_frame_transed_reg[8]_i_1_n_8 ,\good_frame_transed_reg[8]_i_1_n_9 ,\good_frame_transed_reg[8]_i_1_n_10 ,\good_frame_transed_reg[8]_i_1_n_11 ,\good_frame_transed_reg[8]_i_1_n_12 ,\good_frame_transed_reg[8]_i_1_n_13 ,\good_frame_transed_reg[8]_i_1_n_14 ,\good_frame_transed_reg[8]_i_1_n_15 }),
        .S(good_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \good_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[1]),
        .CLR(rst_i),
        .D(\good_frame_transed_reg[8]_i_1_n_14 ),
        .Q(good_frame_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \lt_out_range[0]_i_2 
       (.I0(lt_out_range_reg[0]),
        .O(\lt_out_range[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_15 ),
        .Q(lt_out_range_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[0]_i_1_n_0 ,\lt_out_range_reg[0]_i_1_n_1 ,\lt_out_range_reg[0]_i_1_n_2 ,\lt_out_range_reg[0]_i_1_n_3 ,\lt_out_range_reg[0]_i_1_n_4 ,\lt_out_range_reg[0]_i_1_n_5 ,\lt_out_range_reg[0]_i_1_n_6 ,\lt_out_range_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\lt_out_range_reg[0]_i_1_n_8 ,\lt_out_range_reg[0]_i_1_n_9 ,\lt_out_range_reg[0]_i_1_n_10 ,\lt_out_range_reg[0]_i_1_n_11 ,\lt_out_range_reg[0]_i_1_n_12 ,\lt_out_range_reg[0]_i_1_n_13 ,\lt_out_range_reg[0]_i_1_n_14 ,\lt_out_range_reg[0]_i_1_n_15 }),
        .S({lt_out_range_reg[7:1],\lt_out_range[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_13 ),
        .Q(lt_out_range_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_12 ),
        .Q(lt_out_range_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_11 ),
        .Q(lt_out_range_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_10 ),
        .Q(lt_out_range_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_9 ),
        .Q(lt_out_range_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_8 ),
        .Q(lt_out_range_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_15 ),
        .Q(lt_out_range_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[16]_i_1 
       (.CI(\lt_out_range_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[16]_i_1_n_0 ,\lt_out_range_reg[16]_i_1_n_1 ,\lt_out_range_reg[16]_i_1_n_2 ,\lt_out_range_reg[16]_i_1_n_3 ,\lt_out_range_reg[16]_i_1_n_4 ,\lt_out_range_reg[16]_i_1_n_5 ,\lt_out_range_reg[16]_i_1_n_6 ,\lt_out_range_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[16]_i_1_n_8 ,\lt_out_range_reg[16]_i_1_n_9 ,\lt_out_range_reg[16]_i_1_n_10 ,\lt_out_range_reg[16]_i_1_n_11 ,\lt_out_range_reg[16]_i_1_n_12 ,\lt_out_range_reg[16]_i_1_n_13 ,\lt_out_range_reg[16]_i_1_n_14 ,\lt_out_range_reg[16]_i_1_n_15 }),
        .S(lt_out_range_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_14 ),
        .Q(lt_out_range_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_13 ),
        .Q(lt_out_range_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_12 ),
        .Q(lt_out_range_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_14 ),
        .Q(lt_out_range_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_11 ),
        .Q(lt_out_range_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_10 ),
        .Q(lt_out_range_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_9 ),
        .Q(lt_out_range_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[16]_i_1_n_8 ),
        .Q(lt_out_range_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_15 ),
        .Q(lt_out_range_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[24]_i_1 
       (.CI(\lt_out_range_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[24]_i_1_n_0 ,\lt_out_range_reg[24]_i_1_n_1 ,\lt_out_range_reg[24]_i_1_n_2 ,\lt_out_range_reg[24]_i_1_n_3 ,\lt_out_range_reg[24]_i_1_n_4 ,\lt_out_range_reg[24]_i_1_n_5 ,\lt_out_range_reg[24]_i_1_n_6 ,\lt_out_range_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[24]_i_1_n_8 ,\lt_out_range_reg[24]_i_1_n_9 ,\lt_out_range_reg[24]_i_1_n_10 ,\lt_out_range_reg[24]_i_1_n_11 ,\lt_out_range_reg[24]_i_1_n_12 ,\lt_out_range_reg[24]_i_1_n_13 ,\lt_out_range_reg[24]_i_1_n_14 ,\lt_out_range_reg[24]_i_1_n_15 }),
        .S(lt_out_range_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_14 ),
        .Q(lt_out_range_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_13 ),
        .Q(lt_out_range_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_12 ),
        .Q(lt_out_range_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_11 ),
        .Q(lt_out_range_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_10 ),
        .Q(lt_out_range_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_13 ),
        .Q(lt_out_range_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_9 ),
        .Q(lt_out_range_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[24]_i_1_n_8 ),
        .Q(lt_out_range_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_15 ),
        .Q(lt_out_range_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[32]_i_1 
       (.CI(\lt_out_range_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[32]_i_1_n_0 ,\lt_out_range_reg[32]_i_1_n_1 ,\lt_out_range_reg[32]_i_1_n_2 ,\lt_out_range_reg[32]_i_1_n_3 ,\lt_out_range_reg[32]_i_1_n_4 ,\lt_out_range_reg[32]_i_1_n_5 ,\lt_out_range_reg[32]_i_1_n_6 ,\lt_out_range_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[32]_i_1_n_8 ,\lt_out_range_reg[32]_i_1_n_9 ,\lt_out_range_reg[32]_i_1_n_10 ,\lt_out_range_reg[32]_i_1_n_11 ,\lt_out_range_reg[32]_i_1_n_12 ,\lt_out_range_reg[32]_i_1_n_13 ,\lt_out_range_reg[32]_i_1_n_14 ,\lt_out_range_reg[32]_i_1_n_15 }),
        .S(lt_out_range_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_14 ),
        .Q(lt_out_range_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_13 ),
        .Q(lt_out_range_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_12 ),
        .Q(lt_out_range_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_11 ),
        .Q(lt_out_range_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_10 ),
        .Q(lt_out_range_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_9 ),
        .Q(lt_out_range_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[32]_i_1_n_8 ),
        .Q(lt_out_range_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_12 ),
        .Q(lt_out_range_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_15 ),
        .Q(lt_out_range_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[40]_i_1 
       (.CI(\lt_out_range_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[40]_i_1_n_0 ,\lt_out_range_reg[40]_i_1_n_1 ,\lt_out_range_reg[40]_i_1_n_2 ,\lt_out_range_reg[40]_i_1_n_3 ,\lt_out_range_reg[40]_i_1_n_4 ,\lt_out_range_reg[40]_i_1_n_5 ,\lt_out_range_reg[40]_i_1_n_6 ,\lt_out_range_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[40]_i_1_n_8 ,\lt_out_range_reg[40]_i_1_n_9 ,\lt_out_range_reg[40]_i_1_n_10 ,\lt_out_range_reg[40]_i_1_n_11 ,\lt_out_range_reg[40]_i_1_n_12 ,\lt_out_range_reg[40]_i_1_n_13 ,\lt_out_range_reg[40]_i_1_n_14 ,\lt_out_range_reg[40]_i_1_n_15 }),
        .S(lt_out_range_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_14 ),
        .Q(lt_out_range_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_13 ),
        .Q(lt_out_range_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_12 ),
        .Q(lt_out_range_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_11 ),
        .Q(lt_out_range_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_10 ),
        .Q(lt_out_range_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_9 ),
        .Q(lt_out_range_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[40]_i_1_n_8 ),
        .Q(lt_out_range_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_15 ),
        .Q(lt_out_range_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[48]_i_1 
       (.CI(\lt_out_range_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[48]_i_1_n_0 ,\lt_out_range_reg[48]_i_1_n_1 ,\lt_out_range_reg[48]_i_1_n_2 ,\lt_out_range_reg[48]_i_1_n_3 ,\lt_out_range_reg[48]_i_1_n_4 ,\lt_out_range_reg[48]_i_1_n_5 ,\lt_out_range_reg[48]_i_1_n_6 ,\lt_out_range_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[48]_i_1_n_8 ,\lt_out_range_reg[48]_i_1_n_9 ,\lt_out_range_reg[48]_i_1_n_10 ,\lt_out_range_reg[48]_i_1_n_11 ,\lt_out_range_reg[48]_i_1_n_12 ,\lt_out_range_reg[48]_i_1_n_13 ,\lt_out_range_reg[48]_i_1_n_14 ,\lt_out_range_reg[48]_i_1_n_15 }),
        .S(lt_out_range_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_14 ),
        .Q(lt_out_range_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_11 ),
        .Q(lt_out_range_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_13 ),
        .Q(lt_out_range_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_12 ),
        .Q(lt_out_range_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_11 ),
        .Q(lt_out_range_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_10 ),
        .Q(lt_out_range_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_9 ),
        .Q(lt_out_range_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[48]_i_1_n_8 ),
        .Q(lt_out_range_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_15 ),
        .Q(lt_out_range_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[56]_i_1 
       (.CI(\lt_out_range_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_lt_out_range_reg[56]_i_1_CO_UNCONNECTED [7],\lt_out_range_reg[56]_i_1_n_1 ,\lt_out_range_reg[56]_i_1_n_2 ,\lt_out_range_reg[56]_i_1_n_3 ,\lt_out_range_reg[56]_i_1_n_4 ,\lt_out_range_reg[56]_i_1_n_5 ,\lt_out_range_reg[56]_i_1_n_6 ,\lt_out_range_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[56]_i_1_n_8 ,\lt_out_range_reg[56]_i_1_n_9 ,\lt_out_range_reg[56]_i_1_n_10 ,\lt_out_range_reg[56]_i_1_n_11 ,\lt_out_range_reg[56]_i_1_n_12 ,\lt_out_range_reg[56]_i_1_n_13 ,\lt_out_range_reg[56]_i_1_n_14 ,\lt_out_range_reg[56]_i_1_n_15 }),
        .S(lt_out_range_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_14 ),
        .Q(lt_out_range_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_13 ),
        .Q(lt_out_range_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_12 ),
        .Q(lt_out_range_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_10 ),
        .Q(lt_out_range_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_11 ),
        .Q(lt_out_range_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_10 ),
        .Q(lt_out_range_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_9 ),
        .Q(lt_out_range_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[56]_i_1_n_8 ),
        .Q(lt_out_range_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_9 ),
        .Q(lt_out_range_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[0]_i_1_n_8 ),
        .Q(lt_out_range_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_15 ),
        .Q(lt_out_range_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \lt_out_range_reg[8]_i_1 
       (.CI(\lt_out_range_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\lt_out_range_reg[8]_i_1_n_0 ,\lt_out_range_reg[8]_i_1_n_1 ,\lt_out_range_reg[8]_i_1_n_2 ,\lt_out_range_reg[8]_i_1_n_3 ,\lt_out_range_reg[8]_i_1_n_4 ,\lt_out_range_reg[8]_i_1_n_5 ,\lt_out_range_reg[8]_i_1_n_6 ,\lt_out_range_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\lt_out_range_reg[8]_i_1_n_8 ,\lt_out_range_reg[8]_i_1_n_9 ,\lt_out_range_reg[8]_i_1_n_10 ,\lt_out_range_reg[8]_i_1_n_11 ,\lt_out_range_reg[8]_i_1_n_12 ,\lt_out_range_reg[8]_i_1_n_13 ,\lt_out_range_reg[8]_i_1_n_14 ,\lt_out_range_reg[8]_i_1_n_15 }),
        .S(lt_out_range_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_out_range_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[11]),
        .CLR(rst_i),
        .D(\lt_out_range_reg[8]_i_1_n_14 ),
        .Q(lt_out_range_reg[9]));
  FDCE #(
    .INIT(1'b0)) 
    mdio_in_valid_d1_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(mdio_in_valid),
        .Q(mdio_in_valid_d1));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    \mdio_opcode[1]_i_1 
       (.I0(\recv_config0_reg[0]_0 ),
        .I1(\stat_rd_data_reg[63]_0 ),
        .I2(\stat_rd_data_reg[63]_1 ),
        .I3(mdio_opcode),
        .O(\mdio_opcode[1]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_opcode_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\mdio_opcode[1]_i_1_n_0 ),
        .Q(mdio_opcode));
  LUT4 #(
    .INIT(16'h8F88)) 
    mdio_out_valid_i_1
       (.I0(\stat_rd_data_reg[63]_1 ),
        .I1(\stat_rd_data_reg[63]_0 ),
        .I2(mdio_out_valid_i_2_n_0),
        .I3(mdio_out_valid),
        .O(mdio_out_valid_i_1_n_0));
  LUT5 #(
    .INIT(32'h40000000)) 
    mdio_out_valid_i_2
       (.I0(tmp_cnt[0]),
        .I1(tmp_cnt[1]),
        .I2(tmp_cnt[4]),
        .I3(tmp_cnt[3]),
        .I4(tmp_cnt[2]),
        .O(mdio_out_valid_i_2_n_0));
  FDCE #(
    .INIT(1'b0)) 
    mdio_out_valid_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(mdio_out_valid_i_1_n_0),
        .Q(mdio_out_valid));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_addr_d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(out[4]),
        .Q(sel0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_addr_d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(out[5]),
        .Q(sel0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_addr_d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(out[6]),
        .Q(sel0[2]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_addr_d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(out[7]),
        .Q(sel0[3]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_addr_d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(out[8]),
        .Q(sel0[4]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \mgmt_config[31]_i_1 
       (.I0(recv_config01__0),
        .I1(\recv_config1[31]_i_3_n_0 ),
        .I2(out[7]),
        .I3(out[1]),
        .I4(\mgmt_config[31]_i_2_n_0 ),
        .I5(out[6]),
        .O(\mgmt_config[31]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFFEF)) 
    \mgmt_config[31]_i_2 
       (.I0(out[3]),
        .I1(out[4]),
        .I2(out[8]),
        .I3(out[2]),
        .O(\mgmt_config[31]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[0] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[0]),
        .Q(Q[0]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[10] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[10]),
        .Q(mgmt_config[10]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[11] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[11]),
        .Q(mgmt_config[11]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[12] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[12]),
        .Q(mgmt_config[12]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[13] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[13]),
        .Q(mgmt_config[13]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[14] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[14]),
        .Q(mgmt_config[14]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[15] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[15]),
        .Q(mgmt_config[15]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[16] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[16]),
        .Q(mgmt_config[16]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[17] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[17]),
        .Q(mgmt_config[17]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[18] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[18]),
        .Q(mgmt_config[18]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[19] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[19]),
        .Q(mgmt_config[19]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[1] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[1]),
        .Q(Q[1]));
  FDPE #(
    .INIT(1'b1)) 
    \mgmt_config_reg[20] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .D(mgmt_wr_data[20]),
        .PRE(rst_i),
        .Q(mgmt_config[20]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[21] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[21]),
        .Q(mgmt_config[21]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[22] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[22]),
        .Q(mgmt_config[22]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[23] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[23]),
        .Q(mgmt_config[23]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[24] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[24]),
        .Q(mgmt_config[24]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[25] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[25]),
        .Q(mgmt_config[25]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[26] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[26]),
        .Q(mgmt_config[26]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[27] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[27]),
        .Q(mgmt_config[27]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[28] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[28]),
        .Q(mgmt_config[28]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[29] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[29]),
        .Q(mgmt_config[29]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[2] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[2]),
        .Q(Q[2]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[30] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[30]),
        .Q(mgmt_config[30]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[31] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[31]),
        .Q(mgmt_config[31]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[3] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[3]),
        .Q(Q[3]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[4] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[4]),
        .Q(Q[4]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[5] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[5]),
        .Q(mgmt_config[5]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[6] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[6]),
        .Q(mgmt_config[6]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[7] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[7]),
        .Q(mgmt_config[7]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[8] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[8]),
        .Q(mgmt_config[8]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_config_reg[9] 
       (.C(clk_i),
        .CE(\mgmt_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[9]),
        .Q(mgmt_config[9]));
  LUT6 #(
    .INIT(64'hFFFF305500FF3055)) 
    mgmt_miim_rdy_i_1
       (.I0(state15_out),
        .I1(mdio_in_valid),
        .I2(mdio_in_valid_d1),
        .I3(\state_reg_n_0_[0] ),
        .I4(\state_reg_n_0_[1] ),
        .I5(in0),
        .O(mgmt_miim_rdy_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    mgmt_miim_rdy_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(mgmt_miim_rdy_i_1_n_0),
        .Q(in0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[0]_i_1 
       (.I0(\mgmt_rd_data[0]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[0]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [0]),
        .O(p_1_in[0]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[0]_i_2 
       (.I0(Q[0]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[0] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[0]_i_4_n_0 ),
        .O(\mgmt_rd_data[0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[0]_i_3 
       (.I0(stat_rd_data[32]),
        .I1(data_sel),
        .I2(stat_rd_data[0]),
        .O(mgmt_rd_data0_in[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[0]_i_4 
       (.I0(\flow_control_config_reg_n_0_[0] ),
        .I1(\trans_config_reg_n_0_[0] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[32]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[0]),
        .O(\mgmt_rd_data[0]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[10]_i_1 
       (.I0(\mgmt_rd_data[10]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[10]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [10]),
        .O(p_1_in[10]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[10]_i_2 
       (.I0(mgmt_config[10]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[10] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[10]_i_4_n_0 ),
        .O(\mgmt_rd_data[10]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[10]_i_3 
       (.I0(stat_rd_data[42]),
        .I1(data_sel),
        .I2(stat_rd_data[10]),
        .O(mgmt_rd_data0_in[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[10]_i_4 
       (.I0(\flow_control_config_reg_n_0_[10] ),
        .I1(\trans_config_reg_n_0_[10] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[42]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[10]),
        .O(\mgmt_rd_data[10]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[11]_i_1 
       (.I0(\mgmt_rd_data[11]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[11]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [11]),
        .O(p_1_in[11]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[11]_i_2 
       (.I0(mgmt_config[11]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[11] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[11]_i_4_n_0 ),
        .O(\mgmt_rd_data[11]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[11]_i_3 
       (.I0(stat_rd_data[43]),
        .I1(data_sel),
        .I2(stat_rd_data[11]),
        .O(mgmt_rd_data0_in[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[11]_i_4 
       (.I0(\flow_control_config_reg_n_0_[11] ),
        .I1(\trans_config_reg_n_0_[11] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[43]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[11]),
        .O(\mgmt_rd_data[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[12]_i_1 
       (.I0(\mgmt_rd_data[12]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[12]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [12]),
        .O(p_1_in[12]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[12]_i_2 
       (.I0(mgmt_config[12]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[12] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[12]_i_4_n_0 ),
        .O(\mgmt_rd_data[12]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[12]_i_3 
       (.I0(stat_rd_data[44]),
        .I1(data_sel),
        .I2(stat_rd_data[12]),
        .O(mgmt_rd_data0_in[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[12]_i_4 
       (.I0(\flow_control_config_reg_n_0_[12] ),
        .I1(\trans_config_reg_n_0_[12] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[44]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[12]),
        .O(\mgmt_rd_data[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[13]_i_1 
       (.I0(\mgmt_rd_data[13]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[13]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [13]),
        .O(p_1_in[13]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[13]_i_2 
       (.I0(mgmt_config[13]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[13] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[13]_i_4_n_0 ),
        .O(\mgmt_rd_data[13]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[13]_i_3 
       (.I0(stat_rd_data[45]),
        .I1(data_sel),
        .I2(stat_rd_data[13]),
        .O(mgmt_rd_data0_in[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[13]_i_4 
       (.I0(\flow_control_config_reg_n_0_[13] ),
        .I1(\trans_config_reg_n_0_[13] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[45]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[13]),
        .O(\mgmt_rd_data[13]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[14]_i_1 
       (.I0(\mgmt_rd_data[14]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[14]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [14]),
        .O(p_1_in[14]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[14]_i_2 
       (.I0(mgmt_config[14]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[14] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[14]_i_4_n_0 ),
        .O(\mgmt_rd_data[14]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[14]_i_3 
       (.I0(stat_rd_data[46]),
        .I1(data_sel),
        .I2(stat_rd_data[14]),
        .O(mgmt_rd_data0_in[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[14]_i_4 
       (.I0(\flow_control_config_reg_n_0_[14] ),
        .I1(\trans_config_reg_n_0_[14] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[46]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[14]),
        .O(\mgmt_rd_data[14]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[15]_i_1 
       (.I0(\mgmt_rd_data[15]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[15]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [15]),
        .O(p_1_in[15]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[15]_i_2 
       (.I0(mgmt_config[15]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[15] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[15]_i_4_n_0 ),
        .O(\mgmt_rd_data[15]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[15]_i_3 
       (.I0(stat_rd_data[47]),
        .I1(data_sel),
        .I2(stat_rd_data[15]),
        .O(mgmt_rd_data0_in[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[15]_i_4 
       (.I0(\flow_control_config_reg_n_0_[15] ),
        .I1(\trans_config_reg_n_0_[15] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[47]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[15]),
        .O(\mgmt_rd_data[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[16]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[16]),
        .I2(data_sel),
        .I3(stat_rd_data[48]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[16]_i_2_n_0 ),
        .O(p_1_in[16]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[16]_i_2 
       (.I0(mgmt_config[16]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[16] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[16]_i_3_n_0 ),
        .O(\mgmt_rd_data[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[16]_i_3 
       (.I0(\flow_control_config_reg_n_0_[16] ),
        .I1(\trans_config_reg_n_0_[16] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[16] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[16]),
        .O(\mgmt_rd_data[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[17]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[17]),
        .I2(data_sel),
        .I3(stat_rd_data[49]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[17]_i_2_n_0 ),
        .O(p_1_in[17]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[17]_i_2 
       (.I0(mgmt_config[17]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[17] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[17]_i_3_n_0 ),
        .O(\mgmt_rd_data[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[17]_i_3 
       (.I0(\flow_control_config_reg_n_0_[17] ),
        .I1(\trans_config_reg_n_0_[17] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[17] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[17]),
        .O(\mgmt_rd_data[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[18]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[18]),
        .I2(data_sel),
        .I3(stat_rd_data[50]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[18]_i_2_n_0 ),
        .O(p_1_in[18]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[18]_i_2 
       (.I0(mgmt_config[18]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[18] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[18]_i_3_n_0 ),
        .O(\mgmt_rd_data[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[18]_i_3 
       (.I0(\flow_control_config_reg_n_0_[18] ),
        .I1(\trans_config_reg_n_0_[18] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[18] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[18]),
        .O(\mgmt_rd_data[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[19]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[19]),
        .I2(data_sel),
        .I3(stat_rd_data[51]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[19]_i_2_n_0 ),
        .O(p_1_in[19]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[19]_i_2 
       (.I0(mgmt_config[19]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[19] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[19]_i_3_n_0 ),
        .O(\mgmt_rd_data[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[19]_i_3 
       (.I0(\flow_control_config_reg_n_0_[19] ),
        .I1(\trans_config_reg_n_0_[19] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[19] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[19]),
        .O(\mgmt_rd_data[19]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[1]_i_1 
       (.I0(\mgmt_rd_data[1]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[1]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [1]),
        .O(p_1_in[1]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[1]_i_2 
       (.I0(Q[1]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[1] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[1]_i_4_n_0 ),
        .O(\mgmt_rd_data[1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[1]_i_3 
       (.I0(stat_rd_data[33]),
        .I1(data_sel),
        .I2(stat_rd_data[1]),
        .O(mgmt_rd_data0_in[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[1]_i_4 
       (.I0(\flow_control_config_reg_n_0_[1] ),
        .I1(\trans_config_reg_n_0_[1] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[33]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[1]),
        .O(\mgmt_rd_data[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[20]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[20]),
        .I2(data_sel),
        .I3(stat_rd_data[52]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[20]_i_2_n_0 ),
        .O(p_1_in[20]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[20]_i_2 
       (.I0(mgmt_config[20]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[20] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[20]_i_3_n_0 ),
        .O(\mgmt_rd_data[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[20]_i_3 
       (.I0(\flow_control_config_reg_n_0_[20] ),
        .I1(\trans_config_reg_n_0_[20] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[20] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[20]),
        .O(\mgmt_rd_data[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[21]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[21]),
        .I2(data_sel),
        .I3(stat_rd_data[53]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[21]_i_2_n_0 ),
        .O(p_1_in[21]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[21]_i_2 
       (.I0(mgmt_config[21]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[21] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[21]_i_3_n_0 ),
        .O(\mgmt_rd_data[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[21]_i_3 
       (.I0(\flow_control_config_reg_n_0_[21] ),
        .I1(\trans_config_reg_n_0_[21] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[21] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[21]),
        .O(\mgmt_rd_data[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[22]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[22]),
        .I2(data_sel),
        .I3(stat_rd_data[54]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[22]_i_2_n_0 ),
        .O(p_1_in[22]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[22]_i_2 
       (.I0(mgmt_config[22]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[22] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[22]_i_3_n_0 ),
        .O(\mgmt_rd_data[22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[22]_i_3 
       (.I0(\flow_control_config_reg_n_0_[22] ),
        .I1(\trans_config_reg_n_0_[22] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[22] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[22]),
        .O(\mgmt_rd_data[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[23]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[23]),
        .I2(data_sel),
        .I3(stat_rd_data[55]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[23]_i_2_n_0 ),
        .O(p_1_in[23]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[23]_i_2 
       (.I0(mgmt_config[23]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[23] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[23]_i_3_n_0 ),
        .O(\mgmt_rd_data[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[23]_i_3 
       (.I0(\flow_control_config_reg_n_0_[23] ),
        .I1(\trans_config_reg_n_0_[23] ),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[23] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[23]),
        .O(\mgmt_rd_data[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[24]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[24]),
        .I2(data_sel),
        .I3(stat_rd_data[56]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[24]_i_2_n_0 ),
        .O(p_1_in[24]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[24]_i_2 
       (.I0(mgmt_config[24]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[24] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[24]_i_3_n_0 ),
        .O(\mgmt_rd_data[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[24]_i_3 
       (.I0(\flow_control_config_reg_n_0_[24] ),
        .I1(cfgTxRegData[1]),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[24] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[24]),
        .O(\mgmt_rd_data[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[25]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[25]),
        .I2(data_sel),
        .I3(stat_rd_data[57]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[25]_i_2_n_0 ),
        .O(p_1_in[25]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[25]_i_2 
       (.I0(mgmt_config[25]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[25] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[25]_i_3_n_0 ),
        .O(\mgmt_rd_data[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[25]_i_3 
       (.I0(\flow_control_config_reg_n_0_[25] ),
        .I1(cfgTxRegData[2]),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[25] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[25]),
        .O(\mgmt_rd_data[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[26]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[26]),
        .I2(data_sel),
        .I3(stat_rd_data[58]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[26]_i_2_n_0 ),
        .O(p_1_in[26]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[26]_i_2 
       (.I0(mgmt_config[26]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[26] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[26]_i_3_n_0 ),
        .O(\mgmt_rd_data[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[26]_i_3 
       (.I0(\flow_control_config_reg_n_0_[26] ),
        .I1(cfgTxRegData[3]),
        .I2(sel0[3]),
        .I3(\recv_config1_reg_n_0_[26] ),
        .I4(sel0[2]),
        .I5(cfgRxRegData[26]),
        .O(\mgmt_rd_data[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[27]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[27]),
        .I2(data_sel),
        .I3(stat_rd_data[59]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[27]_i_2_n_0 ),
        .O(p_1_in[27]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[27]_i_2 
       (.I0(mgmt_config[27]),
        .I1(sel0[2]),
        .I2(cfgTxRegData[9]),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[27]_i_3_n_0 ),
        .O(\mgmt_rd_data[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[27]_i_3 
       (.I0(\flow_control_config_reg_n_0_[27] ),
        .I1(cfgTxRegData[4]),
        .I2(sel0[3]),
        .I3(cfgRxRegData[48]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[27]),
        .O(\mgmt_rd_data[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[28]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[28]),
        .I2(data_sel),
        .I3(stat_rd_data[60]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[28]_i_2_n_0 ),
        .O(p_1_in[28]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[28]_i_2 
       (.I0(mgmt_config[28]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[28] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[28]_i_3_n_0 ),
        .O(\mgmt_rd_data[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[28]_i_3 
       (.I0(\flow_control_config_reg_n_0_[28] ),
        .I1(cfgTxRegData[5]),
        .I2(sel0[3]),
        .I3(cfgRxRegData[49]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[28]),
        .O(\mgmt_rd_data[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[29]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[29]),
        .I2(data_sel),
        .I3(stat_rd_data[61]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[29]_i_2_n_0 ),
        .O(p_1_in[29]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[29]_i_2 
       (.I0(mgmt_config[29]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[29] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[29]_i_3_n_0 ),
        .O(\mgmt_rd_data[29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[29]_i_3 
       (.I0(\flow_control_config_reg_n_0_[29] ),
        .I1(cfgTxRegData[6]),
        .I2(sel0[3]),
        .I3(cfgRxRegData[50]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[29]),
        .O(\mgmt_rd_data[29]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[2]_i_1 
       (.I0(\mgmt_rd_data[2]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[2]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [2]),
        .O(p_1_in[2]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[2]_i_2 
       (.I0(Q[2]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[2] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[2]_i_4_n_0 ),
        .O(\mgmt_rd_data[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[2]_i_3 
       (.I0(stat_rd_data[34]),
        .I1(data_sel),
        .I2(stat_rd_data[2]),
        .O(mgmt_rd_data0_in[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[2]_i_4 
       (.I0(\flow_control_config_reg_n_0_[2] ),
        .I1(\trans_config_reg_n_0_[2] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[34]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[2]),
        .O(\mgmt_rd_data[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[30]_i_1 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[30]),
        .I2(data_sel),
        .I3(stat_rd_data[62]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[30]_i_2_n_0 ),
        .O(p_1_in[30]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[30]_i_2 
       (.I0(mgmt_config[30]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[30] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[30]_i_3_n_0 ),
        .O(\mgmt_rd_data[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[30]_i_3 
       (.I0(cfgTxRegData[0]),
        .I1(cfgTxRegData[7]),
        .I2(sel0[3]),
        .I3(cfgRxRegData[51]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[30]),
        .O(\mgmt_rd_data[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h88B88888)) 
    \mgmt_rd_data[31]_i_1 
       (.I0(\mgmt_rd_data[31]_i_3_n_0 ),
        .I1(\state_reg_n_0_[1] ),
        .I2(\state_reg_n_0_[0] ),
        .I3(mdio_in_valid),
        .I4(mdio_in_valid_d1),
        .O(mgmt_rd_data0));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \mgmt_rd_data[31]_i_2 
       (.I0(\state_reg_n_0_[1] ),
        .I1(stat_rd_data[31]),
        .I2(data_sel),
        .I3(stat_rd_data[63]),
        .I4(\state_reg_n_0_[0] ),
        .I5(\mgmt_rd_data[31]_i_4_n_0 ),
        .O(p_1_in[31]));
  LUT5 #(
    .INIT(32'h55575757)) 
    \mgmt_rd_data[31]_i_3 
       (.I0(\state_reg_n_0_[0] ),
        .I1(sel0[1]),
        .I2(sel0[0]),
        .I3(sel0[3]),
        .I4(sel0[4]),
        .O(\mgmt_rd_data[31]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[31]_i_4 
       (.I0(mgmt_config[31]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[31] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[31]_i_5_n_0 ),
        .O(\mgmt_rd_data[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[31]_i_5 
       (.I0(\flow_control_config_reg_n_0_[31] ),
        .I1(cfgTxRegData[8]),
        .I2(sel0[3]),
        .I3(cfgRxRegData[52]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[31]),
        .O(\mgmt_rd_data[31]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[3]_i_1 
       (.I0(\mgmt_rd_data[3]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[3]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [3]),
        .O(p_1_in[3]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[3]_i_2 
       (.I0(Q[3]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[3] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[3]_i_4_n_0 ),
        .O(\mgmt_rd_data[3]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[3]_i_3 
       (.I0(stat_rd_data[35]),
        .I1(data_sel),
        .I2(stat_rd_data[3]),
        .O(mgmt_rd_data0_in[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[3]_i_4 
       (.I0(\flow_control_config_reg_n_0_[3] ),
        .I1(\trans_config_reg_n_0_[3] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[35]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[3]),
        .O(\mgmt_rd_data[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[4]_i_1 
       (.I0(\mgmt_rd_data[4]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[4]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [4]),
        .O(p_1_in[4]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[4]_i_2 
       (.I0(Q[4]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[4] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[4]_i_4_n_0 ),
        .O(\mgmt_rd_data[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[4]_i_3 
       (.I0(stat_rd_data[36]),
        .I1(data_sel),
        .I2(stat_rd_data[4]),
        .O(mgmt_rd_data0_in[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[4]_i_4 
       (.I0(\flow_control_config_reg_n_0_[4] ),
        .I1(\trans_config_reg_n_0_[4] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[36]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[4]),
        .O(\mgmt_rd_data[4]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[5]_i_1 
       (.I0(\mgmt_rd_data[5]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[5]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [5]),
        .O(p_1_in[5]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[5]_i_2 
       (.I0(mgmt_config[5]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[5] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[5]_i_4_n_0 ),
        .O(\mgmt_rd_data[5]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[5]_i_3 
       (.I0(stat_rd_data[37]),
        .I1(data_sel),
        .I2(stat_rd_data[5]),
        .O(mgmt_rd_data0_in[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[5]_i_4 
       (.I0(\flow_control_config_reg_n_0_[5] ),
        .I1(\trans_config_reg_n_0_[5] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[37]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[5]),
        .O(\mgmt_rd_data[5]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[6]_i_1 
       (.I0(\mgmt_rd_data[6]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[6]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [6]),
        .O(p_1_in[6]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[6]_i_2 
       (.I0(mgmt_config[6]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[6] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[6]_i_4_n_0 ),
        .O(\mgmt_rd_data[6]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[6]_i_3 
       (.I0(stat_rd_data[38]),
        .I1(data_sel),
        .I2(stat_rd_data[6]),
        .O(mgmt_rd_data0_in[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[6]_i_4 
       (.I0(\flow_control_config_reg_n_0_[6] ),
        .I1(\trans_config_reg_n_0_[6] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[38]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[6]),
        .O(\mgmt_rd_data[6]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[7]_i_1 
       (.I0(\mgmt_rd_data[7]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[7]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [7]),
        .O(p_1_in[7]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[7]_i_2 
       (.I0(mgmt_config[7]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[7] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[7]_i_4_n_0 ),
        .O(\mgmt_rd_data[7]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[7]_i_3 
       (.I0(stat_rd_data[39]),
        .I1(data_sel),
        .I2(stat_rd_data[7]),
        .O(mgmt_rd_data0_in[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[7]_i_4 
       (.I0(\flow_control_config_reg_n_0_[7] ),
        .I1(\trans_config_reg_n_0_[7] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[39]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[7]),
        .O(\mgmt_rd_data[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[8]_i_1 
       (.I0(\mgmt_rd_data[8]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[8]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [8]),
        .O(p_1_in[8]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[8]_i_2 
       (.I0(mgmt_config[8]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[8] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[8]_i_4_n_0 ),
        .O(\mgmt_rd_data[8]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[8]_i_3 
       (.I0(stat_rd_data[40]),
        .I1(data_sel),
        .I2(stat_rd_data[8]),
        .O(mgmt_rd_data0_in[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[8]_i_4 
       (.I0(\flow_control_config_reg_n_0_[8] ),
        .I1(\trans_config_reg_n_0_[8] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[40]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[8]),
        .O(\mgmt_rd_data[8]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[9]_i_1 
       (.I0(\mgmt_rd_data[9]_i_2_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(mgmt_rd_data0_in[9]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\mgmt_rd_data_reg[15]_0 [9]),
        .O(p_1_in[9]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mgmt_rd_data[9]_i_2 
       (.I0(mgmt_config[9]),
        .I1(sel0[2]),
        .I2(\rs_config_reg_n_0_[9] ),
        .I3(sel0[4]),
        .I4(\mgmt_rd_data[9]_i_4_n_0 ),
        .O(\mgmt_rd_data[9]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mgmt_rd_data[9]_i_3 
       (.I0(stat_rd_data[41]),
        .I1(data_sel),
        .I2(stat_rd_data[9]),
        .O(mgmt_rd_data0_in[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mgmt_rd_data[9]_i_4 
       (.I0(\flow_control_config_reg_n_0_[9] ),
        .I1(\trans_config_reg_n_0_[9] ),
        .I2(sel0[3]),
        .I3(cfgRxRegData[41]),
        .I4(sel0[2]),
        .I5(cfgRxRegData[9]),
        .O(\mgmt_rd_data[9]_i_4_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[0] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[0]),
        .Q(mgmt_rd_data[0]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[10] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[10]),
        .Q(mgmt_rd_data[10]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[11] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[11]),
        .Q(mgmt_rd_data[11]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[12] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[12]),
        .Q(mgmt_rd_data[12]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[13] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[13]),
        .Q(mgmt_rd_data[13]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[14] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[14]),
        .Q(mgmt_rd_data[14]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[15] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[15]),
        .Q(mgmt_rd_data[15]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[16] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[16]),
        .Q(mgmt_rd_data[16]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[17] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[17]),
        .Q(mgmt_rd_data[17]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[18] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[18]),
        .Q(mgmt_rd_data[18]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[19] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[19]),
        .Q(mgmt_rd_data[19]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[1] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[1]),
        .Q(mgmt_rd_data[1]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[20] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[20]),
        .Q(mgmt_rd_data[20]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[21] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[21]),
        .Q(mgmt_rd_data[21]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[22] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[22]),
        .Q(mgmt_rd_data[22]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[23] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[23]),
        .Q(mgmt_rd_data[23]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[24] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[24]),
        .Q(mgmt_rd_data[24]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[25] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[25]),
        .Q(mgmt_rd_data[25]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[26] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[26]),
        .Q(mgmt_rd_data[26]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[27] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[27]),
        .Q(mgmt_rd_data[27]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[28] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[28]),
        .Q(mgmt_rd_data[28]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[29] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[29]),
        .Q(mgmt_rd_data[29]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[2] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[2]),
        .Q(mgmt_rd_data[2]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[30] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[30]),
        .Q(mgmt_rd_data[30]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[31] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[31]),
        .Q(mgmt_rd_data[31]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[3] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[3]),
        .Q(mgmt_rd_data[3]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[4] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[4]),
        .Q(mgmt_rd_data[4]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[5] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[5]),
        .Q(mgmt_rd_data[5]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[6] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[6]),
        .Q(mgmt_rd_data[6]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[7] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[7]),
        .Q(mgmt_rd_data[7]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[8] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[8]),
        .Q(mgmt_rd_data[8]));
  FDCE #(
    .INIT(1'b0)) 
    \mgmt_rd_data_reg[9] 
       (.C(clk_i),
        .CE(mgmt_rd_data0),
        .CLR(rst_i),
        .D(p_1_in[9]),
        .Q(mgmt_rd_data[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \multicast_frame_transed[0]_i_2 
       (.I0(multicast_frame_transed_reg[0]),
        .O(\multicast_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[0]_i_1_n_0 ,\multicast_frame_transed_reg[0]_i_1_n_1 ,\multicast_frame_transed_reg[0]_i_1_n_2 ,\multicast_frame_transed_reg[0]_i_1_n_3 ,\multicast_frame_transed_reg[0]_i_1_n_4 ,\multicast_frame_transed_reg[0]_i_1_n_5 ,\multicast_frame_transed_reg[0]_i_1_n_6 ,\multicast_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\multicast_frame_transed_reg[0]_i_1_n_8 ,\multicast_frame_transed_reg[0]_i_1_n_9 ,\multicast_frame_transed_reg[0]_i_1_n_10 ,\multicast_frame_transed_reg[0]_i_1_n_11 ,\multicast_frame_transed_reg[0]_i_1_n_12 ,\multicast_frame_transed_reg[0]_i_1_n_13 ,\multicast_frame_transed_reg[0]_i_1_n_14 ,\multicast_frame_transed_reg[0]_i_1_n_15 }),
        .S({multicast_frame_transed_reg[7:1],\multicast_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[16]_i_1 
       (.CI(\multicast_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[16]_i_1_n_0 ,\multicast_frame_transed_reg[16]_i_1_n_1 ,\multicast_frame_transed_reg[16]_i_1_n_2 ,\multicast_frame_transed_reg[16]_i_1_n_3 ,\multicast_frame_transed_reg[16]_i_1_n_4 ,\multicast_frame_transed_reg[16]_i_1_n_5 ,\multicast_frame_transed_reg[16]_i_1_n_6 ,\multicast_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[16]_i_1_n_8 ,\multicast_frame_transed_reg[16]_i_1_n_9 ,\multicast_frame_transed_reg[16]_i_1_n_10 ,\multicast_frame_transed_reg[16]_i_1_n_11 ,\multicast_frame_transed_reg[16]_i_1_n_12 ,\multicast_frame_transed_reg[16]_i_1_n_13 ,\multicast_frame_transed_reg[16]_i_1_n_14 ,\multicast_frame_transed_reg[16]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[16]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[24]_i_1 
       (.CI(\multicast_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[24]_i_1_n_0 ,\multicast_frame_transed_reg[24]_i_1_n_1 ,\multicast_frame_transed_reg[24]_i_1_n_2 ,\multicast_frame_transed_reg[24]_i_1_n_3 ,\multicast_frame_transed_reg[24]_i_1_n_4 ,\multicast_frame_transed_reg[24]_i_1_n_5 ,\multicast_frame_transed_reg[24]_i_1_n_6 ,\multicast_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[24]_i_1_n_8 ,\multicast_frame_transed_reg[24]_i_1_n_9 ,\multicast_frame_transed_reg[24]_i_1_n_10 ,\multicast_frame_transed_reg[24]_i_1_n_11 ,\multicast_frame_transed_reg[24]_i_1_n_12 ,\multicast_frame_transed_reg[24]_i_1_n_13 ,\multicast_frame_transed_reg[24]_i_1_n_14 ,\multicast_frame_transed_reg[24]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[24]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[32]_i_1 
       (.CI(\multicast_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[32]_i_1_n_0 ,\multicast_frame_transed_reg[32]_i_1_n_1 ,\multicast_frame_transed_reg[32]_i_1_n_2 ,\multicast_frame_transed_reg[32]_i_1_n_3 ,\multicast_frame_transed_reg[32]_i_1_n_4 ,\multicast_frame_transed_reg[32]_i_1_n_5 ,\multicast_frame_transed_reg[32]_i_1_n_6 ,\multicast_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[32]_i_1_n_8 ,\multicast_frame_transed_reg[32]_i_1_n_9 ,\multicast_frame_transed_reg[32]_i_1_n_10 ,\multicast_frame_transed_reg[32]_i_1_n_11 ,\multicast_frame_transed_reg[32]_i_1_n_12 ,\multicast_frame_transed_reg[32]_i_1_n_13 ,\multicast_frame_transed_reg[32]_i_1_n_14 ,\multicast_frame_transed_reg[32]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[32]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[40]_i_1 
       (.CI(\multicast_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[40]_i_1_n_0 ,\multicast_frame_transed_reg[40]_i_1_n_1 ,\multicast_frame_transed_reg[40]_i_1_n_2 ,\multicast_frame_transed_reg[40]_i_1_n_3 ,\multicast_frame_transed_reg[40]_i_1_n_4 ,\multicast_frame_transed_reg[40]_i_1_n_5 ,\multicast_frame_transed_reg[40]_i_1_n_6 ,\multicast_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[40]_i_1_n_8 ,\multicast_frame_transed_reg[40]_i_1_n_9 ,\multicast_frame_transed_reg[40]_i_1_n_10 ,\multicast_frame_transed_reg[40]_i_1_n_11 ,\multicast_frame_transed_reg[40]_i_1_n_12 ,\multicast_frame_transed_reg[40]_i_1_n_13 ,\multicast_frame_transed_reg[40]_i_1_n_14 ,\multicast_frame_transed_reg[40]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[40]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[48]_i_1 
       (.CI(\multicast_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[48]_i_1_n_0 ,\multicast_frame_transed_reg[48]_i_1_n_1 ,\multicast_frame_transed_reg[48]_i_1_n_2 ,\multicast_frame_transed_reg[48]_i_1_n_3 ,\multicast_frame_transed_reg[48]_i_1_n_4 ,\multicast_frame_transed_reg[48]_i_1_n_5 ,\multicast_frame_transed_reg[48]_i_1_n_6 ,\multicast_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[48]_i_1_n_8 ,\multicast_frame_transed_reg[48]_i_1_n_9 ,\multicast_frame_transed_reg[48]_i_1_n_10 ,\multicast_frame_transed_reg[48]_i_1_n_11 ,\multicast_frame_transed_reg[48]_i_1_n_12 ,\multicast_frame_transed_reg[48]_i_1_n_13 ,\multicast_frame_transed_reg[48]_i_1_n_14 ,\multicast_frame_transed_reg[48]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[48]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[56]_i_1 
       (.CI(\multicast_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_multicast_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\multicast_frame_transed_reg[56]_i_1_n_1 ,\multicast_frame_transed_reg[56]_i_1_n_2 ,\multicast_frame_transed_reg[56]_i_1_n_3 ,\multicast_frame_transed_reg[56]_i_1_n_4 ,\multicast_frame_transed_reg[56]_i_1_n_5 ,\multicast_frame_transed_reg[56]_i_1_n_6 ,\multicast_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[56]_i_1_n_8 ,\multicast_frame_transed_reg[56]_i_1_n_9 ,\multicast_frame_transed_reg[56]_i_1_n_10 ,\multicast_frame_transed_reg[56]_i_1_n_11 ,\multicast_frame_transed_reg[56]_i_1_n_12 ,\multicast_frame_transed_reg[56]_i_1_n_13 ,\multicast_frame_transed_reg[56]_i_1_n_14 ,\multicast_frame_transed_reg[56]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_13 ),
        .Q(multicast_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_12 ),
        .Q(multicast_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_11 ),
        .Q(multicast_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_10 ),
        .Q(multicast_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[56]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_9 ),
        .Q(multicast_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[0]_i_1_n_8 ),
        .Q(multicast_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_15 ),
        .Q(multicast_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_frame_transed_reg[8]_i_1 
       (.CI(\multicast_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_frame_transed_reg[8]_i_1_n_0 ,\multicast_frame_transed_reg[8]_i_1_n_1 ,\multicast_frame_transed_reg[8]_i_1_n_2 ,\multicast_frame_transed_reg[8]_i_1_n_3 ,\multicast_frame_transed_reg[8]_i_1_n_4 ,\multicast_frame_transed_reg[8]_i_1_n_5 ,\multicast_frame_transed_reg[8]_i_1_n_6 ,\multicast_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_frame_transed_reg[8]_i_1_n_8 ,\multicast_frame_transed_reg[8]_i_1_n_9 ,\multicast_frame_transed_reg[8]_i_1_n_10 ,\multicast_frame_transed_reg[8]_i_1_n_11 ,\multicast_frame_transed_reg[8]_i_1_n_12 ,\multicast_frame_transed_reg[8]_i_1_n_13 ,\multicast_frame_transed_reg[8]_i_1_n_14 ,\multicast_frame_transed_reg[8]_i_1_n_15 }),
        .S(multicast_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_frame_transed_reg[8]_i_1_n_14 ),
        .Q(multicast_frame_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \multicast_received_good[0]_i_2 
       (.I0(multicast_received_good_reg[0]),
        .O(\multicast_received_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_15 ),
        .Q(multicast_received_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[0]_i_1_n_0 ,\multicast_received_good_reg[0]_i_1_n_1 ,\multicast_received_good_reg[0]_i_1_n_2 ,\multicast_received_good_reg[0]_i_1_n_3 ,\multicast_received_good_reg[0]_i_1_n_4 ,\multicast_received_good_reg[0]_i_1_n_5 ,\multicast_received_good_reg[0]_i_1_n_6 ,\multicast_received_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\multicast_received_good_reg[0]_i_1_n_8 ,\multicast_received_good_reg[0]_i_1_n_9 ,\multicast_received_good_reg[0]_i_1_n_10 ,\multicast_received_good_reg[0]_i_1_n_11 ,\multicast_received_good_reg[0]_i_1_n_12 ,\multicast_received_good_reg[0]_i_1_n_13 ,\multicast_received_good_reg[0]_i_1_n_14 ,\multicast_received_good_reg[0]_i_1_n_15 }),
        .S({multicast_received_good_reg[7:1],\multicast_received_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_13 ),
        .Q(multicast_received_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_12 ),
        .Q(multicast_received_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_11 ),
        .Q(multicast_received_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_10 ),
        .Q(multicast_received_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_9 ),
        .Q(multicast_received_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_8 ),
        .Q(multicast_received_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_15 ),
        .Q(multicast_received_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[16]_i_1 
       (.CI(\multicast_received_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[16]_i_1_n_0 ,\multicast_received_good_reg[16]_i_1_n_1 ,\multicast_received_good_reg[16]_i_1_n_2 ,\multicast_received_good_reg[16]_i_1_n_3 ,\multicast_received_good_reg[16]_i_1_n_4 ,\multicast_received_good_reg[16]_i_1_n_5 ,\multicast_received_good_reg[16]_i_1_n_6 ,\multicast_received_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[16]_i_1_n_8 ,\multicast_received_good_reg[16]_i_1_n_9 ,\multicast_received_good_reg[16]_i_1_n_10 ,\multicast_received_good_reg[16]_i_1_n_11 ,\multicast_received_good_reg[16]_i_1_n_12 ,\multicast_received_good_reg[16]_i_1_n_13 ,\multicast_received_good_reg[16]_i_1_n_14 ,\multicast_received_good_reg[16]_i_1_n_15 }),
        .S(multicast_received_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_14 ),
        .Q(multicast_received_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_13 ),
        .Q(multicast_received_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_12 ),
        .Q(multicast_received_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_14 ),
        .Q(multicast_received_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_11 ),
        .Q(multicast_received_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_10 ),
        .Q(multicast_received_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_9 ),
        .Q(multicast_received_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[16]_i_1_n_8 ),
        .Q(multicast_received_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_15 ),
        .Q(multicast_received_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[24]_i_1 
       (.CI(\multicast_received_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[24]_i_1_n_0 ,\multicast_received_good_reg[24]_i_1_n_1 ,\multicast_received_good_reg[24]_i_1_n_2 ,\multicast_received_good_reg[24]_i_1_n_3 ,\multicast_received_good_reg[24]_i_1_n_4 ,\multicast_received_good_reg[24]_i_1_n_5 ,\multicast_received_good_reg[24]_i_1_n_6 ,\multicast_received_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[24]_i_1_n_8 ,\multicast_received_good_reg[24]_i_1_n_9 ,\multicast_received_good_reg[24]_i_1_n_10 ,\multicast_received_good_reg[24]_i_1_n_11 ,\multicast_received_good_reg[24]_i_1_n_12 ,\multicast_received_good_reg[24]_i_1_n_13 ,\multicast_received_good_reg[24]_i_1_n_14 ,\multicast_received_good_reg[24]_i_1_n_15 }),
        .S(multicast_received_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_14 ),
        .Q(multicast_received_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_13 ),
        .Q(multicast_received_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_12 ),
        .Q(multicast_received_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_11 ),
        .Q(multicast_received_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_10 ),
        .Q(multicast_received_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_13 ),
        .Q(multicast_received_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_9 ),
        .Q(multicast_received_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[24]_i_1_n_8 ),
        .Q(multicast_received_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_15 ),
        .Q(multicast_received_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[32]_i_1 
       (.CI(\multicast_received_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[32]_i_1_n_0 ,\multicast_received_good_reg[32]_i_1_n_1 ,\multicast_received_good_reg[32]_i_1_n_2 ,\multicast_received_good_reg[32]_i_1_n_3 ,\multicast_received_good_reg[32]_i_1_n_4 ,\multicast_received_good_reg[32]_i_1_n_5 ,\multicast_received_good_reg[32]_i_1_n_6 ,\multicast_received_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[32]_i_1_n_8 ,\multicast_received_good_reg[32]_i_1_n_9 ,\multicast_received_good_reg[32]_i_1_n_10 ,\multicast_received_good_reg[32]_i_1_n_11 ,\multicast_received_good_reg[32]_i_1_n_12 ,\multicast_received_good_reg[32]_i_1_n_13 ,\multicast_received_good_reg[32]_i_1_n_14 ,\multicast_received_good_reg[32]_i_1_n_15 }),
        .S(multicast_received_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_14 ),
        .Q(multicast_received_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_13 ),
        .Q(multicast_received_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_12 ),
        .Q(multicast_received_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_11 ),
        .Q(multicast_received_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_10 ),
        .Q(multicast_received_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_9 ),
        .Q(multicast_received_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[32]_i_1_n_8 ),
        .Q(multicast_received_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_12 ),
        .Q(multicast_received_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_15 ),
        .Q(multicast_received_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[40]_i_1 
       (.CI(\multicast_received_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[40]_i_1_n_0 ,\multicast_received_good_reg[40]_i_1_n_1 ,\multicast_received_good_reg[40]_i_1_n_2 ,\multicast_received_good_reg[40]_i_1_n_3 ,\multicast_received_good_reg[40]_i_1_n_4 ,\multicast_received_good_reg[40]_i_1_n_5 ,\multicast_received_good_reg[40]_i_1_n_6 ,\multicast_received_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[40]_i_1_n_8 ,\multicast_received_good_reg[40]_i_1_n_9 ,\multicast_received_good_reg[40]_i_1_n_10 ,\multicast_received_good_reg[40]_i_1_n_11 ,\multicast_received_good_reg[40]_i_1_n_12 ,\multicast_received_good_reg[40]_i_1_n_13 ,\multicast_received_good_reg[40]_i_1_n_14 ,\multicast_received_good_reg[40]_i_1_n_15 }),
        .S(multicast_received_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_14 ),
        .Q(multicast_received_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_13 ),
        .Q(multicast_received_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_12 ),
        .Q(multicast_received_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_11 ),
        .Q(multicast_received_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_10 ),
        .Q(multicast_received_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_9 ),
        .Q(multicast_received_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[40]_i_1_n_8 ),
        .Q(multicast_received_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_15 ),
        .Q(multicast_received_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[48]_i_1 
       (.CI(\multicast_received_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[48]_i_1_n_0 ,\multicast_received_good_reg[48]_i_1_n_1 ,\multicast_received_good_reg[48]_i_1_n_2 ,\multicast_received_good_reg[48]_i_1_n_3 ,\multicast_received_good_reg[48]_i_1_n_4 ,\multicast_received_good_reg[48]_i_1_n_5 ,\multicast_received_good_reg[48]_i_1_n_6 ,\multicast_received_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[48]_i_1_n_8 ,\multicast_received_good_reg[48]_i_1_n_9 ,\multicast_received_good_reg[48]_i_1_n_10 ,\multicast_received_good_reg[48]_i_1_n_11 ,\multicast_received_good_reg[48]_i_1_n_12 ,\multicast_received_good_reg[48]_i_1_n_13 ,\multicast_received_good_reg[48]_i_1_n_14 ,\multicast_received_good_reg[48]_i_1_n_15 }),
        .S(multicast_received_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_14 ),
        .Q(multicast_received_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_11 ),
        .Q(multicast_received_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_13 ),
        .Q(multicast_received_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_12 ),
        .Q(multicast_received_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_11 ),
        .Q(multicast_received_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_10 ),
        .Q(multicast_received_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_9 ),
        .Q(multicast_received_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[48]_i_1_n_8 ),
        .Q(multicast_received_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_15 ),
        .Q(multicast_received_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[56]_i_1 
       (.CI(\multicast_received_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_multicast_received_good_reg[56]_i_1_CO_UNCONNECTED [7],\multicast_received_good_reg[56]_i_1_n_1 ,\multicast_received_good_reg[56]_i_1_n_2 ,\multicast_received_good_reg[56]_i_1_n_3 ,\multicast_received_good_reg[56]_i_1_n_4 ,\multicast_received_good_reg[56]_i_1_n_5 ,\multicast_received_good_reg[56]_i_1_n_6 ,\multicast_received_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[56]_i_1_n_8 ,\multicast_received_good_reg[56]_i_1_n_9 ,\multicast_received_good_reg[56]_i_1_n_10 ,\multicast_received_good_reg[56]_i_1_n_11 ,\multicast_received_good_reg[56]_i_1_n_12 ,\multicast_received_good_reg[56]_i_1_n_13 ,\multicast_received_good_reg[56]_i_1_n_14 ,\multicast_received_good_reg[56]_i_1_n_15 }),
        .S(multicast_received_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_14 ),
        .Q(multicast_received_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_13 ),
        .Q(multicast_received_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_12 ),
        .Q(multicast_received_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_10 ),
        .Q(multicast_received_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_11 ),
        .Q(multicast_received_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_10 ),
        .Q(multicast_received_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_9 ),
        .Q(multicast_received_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[56]_i_1_n_8 ),
        .Q(multicast_received_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_9 ),
        .Q(multicast_received_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[0]_i_1_n_8 ),
        .Q(multicast_received_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_15 ),
        .Q(multicast_received_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \multicast_received_good_reg[8]_i_1 
       (.CI(\multicast_received_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\multicast_received_good_reg[8]_i_1_n_0 ,\multicast_received_good_reg[8]_i_1_n_1 ,\multicast_received_good_reg[8]_i_1_n_2 ,\multicast_received_good_reg[8]_i_1_n_3 ,\multicast_received_good_reg[8]_i_1_n_4 ,\multicast_received_good_reg[8]_i_1_n_5 ,\multicast_received_good_reg[8]_i_1_n_6 ,\multicast_received_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\multicast_received_good_reg[8]_i_1_n_8 ,\multicast_received_good_reg[8]_i_1_n_9 ,\multicast_received_good_reg[8]_i_1_n_10 ,\multicast_received_good_reg[8]_i_1_n_11 ,\multicast_received_good_reg[8]_i_1_n_12 ,\multicast_received_good_reg[8]_i_1_n_13 ,\multicast_received_good_reg[8]_i_1_n_14 ,\multicast_received_good_reg[8]_i_1_n_15 }),
        .S(multicast_received_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \multicast_received_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[3]),
        .CLR(rst_i),
        .D(\multicast_received_good_reg[8]_i_1_n_14 ),
        .Q(multicast_received_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \oversize_frame_good[0]_i_2 
       (.I0(oversize_frame_good_reg[0]),
        .O(\oversize_frame_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[0]_i_1_n_0 ,\oversize_frame_good_reg[0]_i_1_n_1 ,\oversize_frame_good_reg[0]_i_1_n_2 ,\oversize_frame_good_reg[0]_i_1_n_3 ,\oversize_frame_good_reg[0]_i_1_n_4 ,\oversize_frame_good_reg[0]_i_1_n_5 ,\oversize_frame_good_reg[0]_i_1_n_6 ,\oversize_frame_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\oversize_frame_good_reg[0]_i_1_n_8 ,\oversize_frame_good_reg[0]_i_1_n_9 ,\oversize_frame_good_reg[0]_i_1_n_10 ,\oversize_frame_good_reg[0]_i_1_n_11 ,\oversize_frame_good_reg[0]_i_1_n_12 ,\oversize_frame_good_reg[0]_i_1_n_13 ,\oversize_frame_good_reg[0]_i_1_n_14 ,\oversize_frame_good_reg[0]_i_1_n_15 }),
        .S({oversize_frame_good_reg[7:1],\oversize_frame_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[16]_i_1 
       (.CI(\oversize_frame_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[16]_i_1_n_0 ,\oversize_frame_good_reg[16]_i_1_n_1 ,\oversize_frame_good_reg[16]_i_1_n_2 ,\oversize_frame_good_reg[16]_i_1_n_3 ,\oversize_frame_good_reg[16]_i_1_n_4 ,\oversize_frame_good_reg[16]_i_1_n_5 ,\oversize_frame_good_reg[16]_i_1_n_6 ,\oversize_frame_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[16]_i_1_n_8 ,\oversize_frame_good_reg[16]_i_1_n_9 ,\oversize_frame_good_reg[16]_i_1_n_10 ,\oversize_frame_good_reg[16]_i_1_n_11 ,\oversize_frame_good_reg[16]_i_1_n_12 ,\oversize_frame_good_reg[16]_i_1_n_13 ,\oversize_frame_good_reg[16]_i_1_n_14 ,\oversize_frame_good_reg[16]_i_1_n_15 }),
        .S(oversize_frame_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[16]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[24]_i_1 
       (.CI(\oversize_frame_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[24]_i_1_n_0 ,\oversize_frame_good_reg[24]_i_1_n_1 ,\oversize_frame_good_reg[24]_i_1_n_2 ,\oversize_frame_good_reg[24]_i_1_n_3 ,\oversize_frame_good_reg[24]_i_1_n_4 ,\oversize_frame_good_reg[24]_i_1_n_5 ,\oversize_frame_good_reg[24]_i_1_n_6 ,\oversize_frame_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[24]_i_1_n_8 ,\oversize_frame_good_reg[24]_i_1_n_9 ,\oversize_frame_good_reg[24]_i_1_n_10 ,\oversize_frame_good_reg[24]_i_1_n_11 ,\oversize_frame_good_reg[24]_i_1_n_12 ,\oversize_frame_good_reg[24]_i_1_n_13 ,\oversize_frame_good_reg[24]_i_1_n_14 ,\oversize_frame_good_reg[24]_i_1_n_15 }),
        .S(oversize_frame_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[24]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[32]_i_1 
       (.CI(\oversize_frame_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[32]_i_1_n_0 ,\oversize_frame_good_reg[32]_i_1_n_1 ,\oversize_frame_good_reg[32]_i_1_n_2 ,\oversize_frame_good_reg[32]_i_1_n_3 ,\oversize_frame_good_reg[32]_i_1_n_4 ,\oversize_frame_good_reg[32]_i_1_n_5 ,\oversize_frame_good_reg[32]_i_1_n_6 ,\oversize_frame_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[32]_i_1_n_8 ,\oversize_frame_good_reg[32]_i_1_n_9 ,\oversize_frame_good_reg[32]_i_1_n_10 ,\oversize_frame_good_reg[32]_i_1_n_11 ,\oversize_frame_good_reg[32]_i_1_n_12 ,\oversize_frame_good_reg[32]_i_1_n_13 ,\oversize_frame_good_reg[32]_i_1_n_14 ,\oversize_frame_good_reg[32]_i_1_n_15 }),
        .S(oversize_frame_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[32]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[40]_i_1 
       (.CI(\oversize_frame_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[40]_i_1_n_0 ,\oversize_frame_good_reg[40]_i_1_n_1 ,\oversize_frame_good_reg[40]_i_1_n_2 ,\oversize_frame_good_reg[40]_i_1_n_3 ,\oversize_frame_good_reg[40]_i_1_n_4 ,\oversize_frame_good_reg[40]_i_1_n_5 ,\oversize_frame_good_reg[40]_i_1_n_6 ,\oversize_frame_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[40]_i_1_n_8 ,\oversize_frame_good_reg[40]_i_1_n_9 ,\oversize_frame_good_reg[40]_i_1_n_10 ,\oversize_frame_good_reg[40]_i_1_n_11 ,\oversize_frame_good_reg[40]_i_1_n_12 ,\oversize_frame_good_reg[40]_i_1_n_13 ,\oversize_frame_good_reg[40]_i_1_n_14 ,\oversize_frame_good_reg[40]_i_1_n_15 }),
        .S(oversize_frame_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[40]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[48]_i_1 
       (.CI(\oversize_frame_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[48]_i_1_n_0 ,\oversize_frame_good_reg[48]_i_1_n_1 ,\oversize_frame_good_reg[48]_i_1_n_2 ,\oversize_frame_good_reg[48]_i_1_n_3 ,\oversize_frame_good_reg[48]_i_1_n_4 ,\oversize_frame_good_reg[48]_i_1_n_5 ,\oversize_frame_good_reg[48]_i_1_n_6 ,\oversize_frame_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[48]_i_1_n_8 ,\oversize_frame_good_reg[48]_i_1_n_9 ,\oversize_frame_good_reg[48]_i_1_n_10 ,\oversize_frame_good_reg[48]_i_1_n_11 ,\oversize_frame_good_reg[48]_i_1_n_12 ,\oversize_frame_good_reg[48]_i_1_n_13 ,\oversize_frame_good_reg[48]_i_1_n_14 ,\oversize_frame_good_reg[48]_i_1_n_15 }),
        .S(oversize_frame_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[48]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[56]_i_1 
       (.CI(\oversize_frame_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_oversize_frame_good_reg[56]_i_1_CO_UNCONNECTED [7],\oversize_frame_good_reg[56]_i_1_n_1 ,\oversize_frame_good_reg[56]_i_1_n_2 ,\oversize_frame_good_reg[56]_i_1_n_3 ,\oversize_frame_good_reg[56]_i_1_n_4 ,\oversize_frame_good_reg[56]_i_1_n_5 ,\oversize_frame_good_reg[56]_i_1_n_6 ,\oversize_frame_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[56]_i_1_n_8 ,\oversize_frame_good_reg[56]_i_1_n_9 ,\oversize_frame_good_reg[56]_i_1_n_10 ,\oversize_frame_good_reg[56]_i_1_n_11 ,\oversize_frame_good_reg[56]_i_1_n_12 ,\oversize_frame_good_reg[56]_i_1_n_13 ,\oversize_frame_good_reg[56]_i_1_n_14 ,\oversize_frame_good_reg[56]_i_1_n_15 }),
        .S(oversize_frame_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_13 ),
        .Q(oversize_frame_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_12 ),
        .Q(oversize_frame_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_11 ),
        .Q(oversize_frame_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_10 ),
        .Q(oversize_frame_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[56]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_9 ),
        .Q(oversize_frame_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[0]_i_1_n_8 ),
        .Q(oversize_frame_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_15 ),
        .Q(oversize_frame_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_good_reg[8]_i_1 
       (.CI(\oversize_frame_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_good_reg[8]_i_1_n_0 ,\oversize_frame_good_reg[8]_i_1_n_1 ,\oversize_frame_good_reg[8]_i_1_n_2 ,\oversize_frame_good_reg[8]_i_1_n_3 ,\oversize_frame_good_reg[8]_i_1_n_4 ,\oversize_frame_good_reg[8]_i_1_n_5 ,\oversize_frame_good_reg[8]_i_1_n_6 ,\oversize_frame_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_good_reg[8]_i_1_n_8 ,\oversize_frame_good_reg[8]_i_1_n_9 ,\oversize_frame_good_reg[8]_i_1_n_10 ,\oversize_frame_good_reg[8]_i_1_n_11 ,\oversize_frame_good_reg[8]_i_1_n_12 ,\oversize_frame_good_reg[8]_i_1_n_13 ,\oversize_frame_good_reg[8]_i_1_n_14 ,\oversize_frame_good_reg[8]_i_1_n_15 }),
        .S(oversize_frame_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[15]),
        .CLR(rst_i),
        .D(\oversize_frame_good_reg[8]_i_1_n_14 ),
        .Q(oversize_frame_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \oversize_frame_transed[0]_i_2 
       (.I0(oversize_frame_transed_reg[0]),
        .O(\oversize_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[0]_i_1_n_0 ,\oversize_frame_transed_reg[0]_i_1_n_1 ,\oversize_frame_transed_reg[0]_i_1_n_2 ,\oversize_frame_transed_reg[0]_i_1_n_3 ,\oversize_frame_transed_reg[0]_i_1_n_4 ,\oversize_frame_transed_reg[0]_i_1_n_5 ,\oversize_frame_transed_reg[0]_i_1_n_6 ,\oversize_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\oversize_frame_transed_reg[0]_i_1_n_8 ,\oversize_frame_transed_reg[0]_i_1_n_9 ,\oversize_frame_transed_reg[0]_i_1_n_10 ,\oversize_frame_transed_reg[0]_i_1_n_11 ,\oversize_frame_transed_reg[0]_i_1_n_12 ,\oversize_frame_transed_reg[0]_i_1_n_13 ,\oversize_frame_transed_reg[0]_i_1_n_14 ,\oversize_frame_transed_reg[0]_i_1_n_15 }),
        .S({oversize_frame_transed_reg[7:1],\oversize_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[16]_i_1 
       (.CI(\oversize_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[16]_i_1_n_0 ,\oversize_frame_transed_reg[16]_i_1_n_1 ,\oversize_frame_transed_reg[16]_i_1_n_2 ,\oversize_frame_transed_reg[16]_i_1_n_3 ,\oversize_frame_transed_reg[16]_i_1_n_4 ,\oversize_frame_transed_reg[16]_i_1_n_5 ,\oversize_frame_transed_reg[16]_i_1_n_6 ,\oversize_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[16]_i_1_n_8 ,\oversize_frame_transed_reg[16]_i_1_n_9 ,\oversize_frame_transed_reg[16]_i_1_n_10 ,\oversize_frame_transed_reg[16]_i_1_n_11 ,\oversize_frame_transed_reg[16]_i_1_n_12 ,\oversize_frame_transed_reg[16]_i_1_n_13 ,\oversize_frame_transed_reg[16]_i_1_n_14 ,\oversize_frame_transed_reg[16]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[16]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[24]_i_1 
       (.CI(\oversize_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[24]_i_1_n_0 ,\oversize_frame_transed_reg[24]_i_1_n_1 ,\oversize_frame_transed_reg[24]_i_1_n_2 ,\oversize_frame_transed_reg[24]_i_1_n_3 ,\oversize_frame_transed_reg[24]_i_1_n_4 ,\oversize_frame_transed_reg[24]_i_1_n_5 ,\oversize_frame_transed_reg[24]_i_1_n_6 ,\oversize_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[24]_i_1_n_8 ,\oversize_frame_transed_reg[24]_i_1_n_9 ,\oversize_frame_transed_reg[24]_i_1_n_10 ,\oversize_frame_transed_reg[24]_i_1_n_11 ,\oversize_frame_transed_reg[24]_i_1_n_12 ,\oversize_frame_transed_reg[24]_i_1_n_13 ,\oversize_frame_transed_reg[24]_i_1_n_14 ,\oversize_frame_transed_reg[24]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[24]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[32]_i_1 
       (.CI(\oversize_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[32]_i_1_n_0 ,\oversize_frame_transed_reg[32]_i_1_n_1 ,\oversize_frame_transed_reg[32]_i_1_n_2 ,\oversize_frame_transed_reg[32]_i_1_n_3 ,\oversize_frame_transed_reg[32]_i_1_n_4 ,\oversize_frame_transed_reg[32]_i_1_n_5 ,\oversize_frame_transed_reg[32]_i_1_n_6 ,\oversize_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[32]_i_1_n_8 ,\oversize_frame_transed_reg[32]_i_1_n_9 ,\oversize_frame_transed_reg[32]_i_1_n_10 ,\oversize_frame_transed_reg[32]_i_1_n_11 ,\oversize_frame_transed_reg[32]_i_1_n_12 ,\oversize_frame_transed_reg[32]_i_1_n_13 ,\oversize_frame_transed_reg[32]_i_1_n_14 ,\oversize_frame_transed_reg[32]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[32]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[40]_i_1 
       (.CI(\oversize_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[40]_i_1_n_0 ,\oversize_frame_transed_reg[40]_i_1_n_1 ,\oversize_frame_transed_reg[40]_i_1_n_2 ,\oversize_frame_transed_reg[40]_i_1_n_3 ,\oversize_frame_transed_reg[40]_i_1_n_4 ,\oversize_frame_transed_reg[40]_i_1_n_5 ,\oversize_frame_transed_reg[40]_i_1_n_6 ,\oversize_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[40]_i_1_n_8 ,\oversize_frame_transed_reg[40]_i_1_n_9 ,\oversize_frame_transed_reg[40]_i_1_n_10 ,\oversize_frame_transed_reg[40]_i_1_n_11 ,\oversize_frame_transed_reg[40]_i_1_n_12 ,\oversize_frame_transed_reg[40]_i_1_n_13 ,\oversize_frame_transed_reg[40]_i_1_n_14 ,\oversize_frame_transed_reg[40]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[40]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[48]_i_1 
       (.CI(\oversize_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[48]_i_1_n_0 ,\oversize_frame_transed_reg[48]_i_1_n_1 ,\oversize_frame_transed_reg[48]_i_1_n_2 ,\oversize_frame_transed_reg[48]_i_1_n_3 ,\oversize_frame_transed_reg[48]_i_1_n_4 ,\oversize_frame_transed_reg[48]_i_1_n_5 ,\oversize_frame_transed_reg[48]_i_1_n_6 ,\oversize_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[48]_i_1_n_8 ,\oversize_frame_transed_reg[48]_i_1_n_9 ,\oversize_frame_transed_reg[48]_i_1_n_10 ,\oversize_frame_transed_reg[48]_i_1_n_11 ,\oversize_frame_transed_reg[48]_i_1_n_12 ,\oversize_frame_transed_reg[48]_i_1_n_13 ,\oversize_frame_transed_reg[48]_i_1_n_14 ,\oversize_frame_transed_reg[48]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[48]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[56]_i_1 
       (.CI(\oversize_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_oversize_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\oversize_frame_transed_reg[56]_i_1_n_1 ,\oversize_frame_transed_reg[56]_i_1_n_2 ,\oversize_frame_transed_reg[56]_i_1_n_3 ,\oversize_frame_transed_reg[56]_i_1_n_4 ,\oversize_frame_transed_reg[56]_i_1_n_5 ,\oversize_frame_transed_reg[56]_i_1_n_6 ,\oversize_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[56]_i_1_n_8 ,\oversize_frame_transed_reg[56]_i_1_n_9 ,\oversize_frame_transed_reg[56]_i_1_n_10 ,\oversize_frame_transed_reg[56]_i_1_n_11 ,\oversize_frame_transed_reg[56]_i_1_n_12 ,\oversize_frame_transed_reg[56]_i_1_n_13 ,\oversize_frame_transed_reg[56]_i_1_n_14 ,\oversize_frame_transed_reg[56]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_13 ),
        .Q(oversize_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_12 ),
        .Q(oversize_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_11 ),
        .Q(oversize_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_10 ),
        .Q(oversize_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[56]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_9 ),
        .Q(oversize_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[0]_i_1_n_8 ),
        .Q(oversize_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_15 ),
        .Q(oversize_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \oversize_frame_transed_reg[8]_i_1 
       (.CI(\oversize_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\oversize_frame_transed_reg[8]_i_1_n_0 ,\oversize_frame_transed_reg[8]_i_1_n_1 ,\oversize_frame_transed_reg[8]_i_1_n_2 ,\oversize_frame_transed_reg[8]_i_1_n_3 ,\oversize_frame_transed_reg[8]_i_1_n_4 ,\oversize_frame_transed_reg[8]_i_1_n_5 ,\oversize_frame_transed_reg[8]_i_1_n_6 ,\oversize_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\oversize_frame_transed_reg[8]_i_1_n_8 ,\oversize_frame_transed_reg[8]_i_1_n_9 ,\oversize_frame_transed_reg[8]_i_1_n_10 ,\oversize_frame_transed_reg[8]_i_1_n_11 ,\oversize_frame_transed_reg[8]_i_1_n_12 ,\oversize_frame_transed_reg[8]_i_1_n_13 ,\oversize_frame_transed_reg[8]_i_1_n_14 ,\oversize_frame_transed_reg[8]_i_1_n_15 }),
        .S(oversize_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \oversize_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[14]),
        .CLR(rst_i),
        .D(\oversize_frame_transed_reg[8]_i_1_n_14 ),
        .Q(oversize_frame_transed_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \pause_frame_good[0]_i_2 
       (.I0(pause_frame_good_reg[0]),
        .O(\pause_frame_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_15 ),
        .Q(pause_frame_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[0]_i_1_n_0 ,\pause_frame_good_reg[0]_i_1_n_1 ,\pause_frame_good_reg[0]_i_1_n_2 ,\pause_frame_good_reg[0]_i_1_n_3 ,\pause_frame_good_reg[0]_i_1_n_4 ,\pause_frame_good_reg[0]_i_1_n_5 ,\pause_frame_good_reg[0]_i_1_n_6 ,\pause_frame_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\pause_frame_good_reg[0]_i_1_n_8 ,\pause_frame_good_reg[0]_i_1_n_9 ,\pause_frame_good_reg[0]_i_1_n_10 ,\pause_frame_good_reg[0]_i_1_n_11 ,\pause_frame_good_reg[0]_i_1_n_12 ,\pause_frame_good_reg[0]_i_1_n_13 ,\pause_frame_good_reg[0]_i_1_n_14 ,\pause_frame_good_reg[0]_i_1_n_15 }),
        .S({pause_frame_good_reg[7:1],\pause_frame_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_13 ),
        .Q(pause_frame_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_12 ),
        .Q(pause_frame_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_11 ),
        .Q(pause_frame_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_10 ),
        .Q(pause_frame_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_9 ),
        .Q(pause_frame_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_8 ),
        .Q(pause_frame_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_15 ),
        .Q(pause_frame_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[16]_i_1 
       (.CI(\pause_frame_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[16]_i_1_n_0 ,\pause_frame_good_reg[16]_i_1_n_1 ,\pause_frame_good_reg[16]_i_1_n_2 ,\pause_frame_good_reg[16]_i_1_n_3 ,\pause_frame_good_reg[16]_i_1_n_4 ,\pause_frame_good_reg[16]_i_1_n_5 ,\pause_frame_good_reg[16]_i_1_n_6 ,\pause_frame_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[16]_i_1_n_8 ,\pause_frame_good_reg[16]_i_1_n_9 ,\pause_frame_good_reg[16]_i_1_n_10 ,\pause_frame_good_reg[16]_i_1_n_11 ,\pause_frame_good_reg[16]_i_1_n_12 ,\pause_frame_good_reg[16]_i_1_n_13 ,\pause_frame_good_reg[16]_i_1_n_14 ,\pause_frame_good_reg[16]_i_1_n_15 }),
        .S(pause_frame_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_14 ),
        .Q(pause_frame_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_13 ),
        .Q(pause_frame_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_12 ),
        .Q(pause_frame_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_14 ),
        .Q(pause_frame_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_11 ),
        .Q(pause_frame_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_10 ),
        .Q(pause_frame_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_9 ),
        .Q(pause_frame_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[16]_i_1_n_8 ),
        .Q(pause_frame_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_15 ),
        .Q(pause_frame_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[24]_i_1 
       (.CI(\pause_frame_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[24]_i_1_n_0 ,\pause_frame_good_reg[24]_i_1_n_1 ,\pause_frame_good_reg[24]_i_1_n_2 ,\pause_frame_good_reg[24]_i_1_n_3 ,\pause_frame_good_reg[24]_i_1_n_4 ,\pause_frame_good_reg[24]_i_1_n_5 ,\pause_frame_good_reg[24]_i_1_n_6 ,\pause_frame_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[24]_i_1_n_8 ,\pause_frame_good_reg[24]_i_1_n_9 ,\pause_frame_good_reg[24]_i_1_n_10 ,\pause_frame_good_reg[24]_i_1_n_11 ,\pause_frame_good_reg[24]_i_1_n_12 ,\pause_frame_good_reg[24]_i_1_n_13 ,\pause_frame_good_reg[24]_i_1_n_14 ,\pause_frame_good_reg[24]_i_1_n_15 }),
        .S(pause_frame_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_14 ),
        .Q(pause_frame_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_13 ),
        .Q(pause_frame_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_12 ),
        .Q(pause_frame_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_11 ),
        .Q(pause_frame_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_10 ),
        .Q(pause_frame_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_13 ),
        .Q(pause_frame_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_9 ),
        .Q(pause_frame_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[24]_i_1_n_8 ),
        .Q(pause_frame_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_15 ),
        .Q(pause_frame_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[32]_i_1 
       (.CI(\pause_frame_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[32]_i_1_n_0 ,\pause_frame_good_reg[32]_i_1_n_1 ,\pause_frame_good_reg[32]_i_1_n_2 ,\pause_frame_good_reg[32]_i_1_n_3 ,\pause_frame_good_reg[32]_i_1_n_4 ,\pause_frame_good_reg[32]_i_1_n_5 ,\pause_frame_good_reg[32]_i_1_n_6 ,\pause_frame_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[32]_i_1_n_8 ,\pause_frame_good_reg[32]_i_1_n_9 ,\pause_frame_good_reg[32]_i_1_n_10 ,\pause_frame_good_reg[32]_i_1_n_11 ,\pause_frame_good_reg[32]_i_1_n_12 ,\pause_frame_good_reg[32]_i_1_n_13 ,\pause_frame_good_reg[32]_i_1_n_14 ,\pause_frame_good_reg[32]_i_1_n_15 }),
        .S(pause_frame_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_14 ),
        .Q(pause_frame_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_13 ),
        .Q(pause_frame_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_12 ),
        .Q(pause_frame_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_11 ),
        .Q(pause_frame_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_10 ),
        .Q(pause_frame_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_9 ),
        .Q(pause_frame_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[32]_i_1_n_8 ),
        .Q(pause_frame_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_12 ),
        .Q(pause_frame_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_15 ),
        .Q(pause_frame_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[40]_i_1 
       (.CI(\pause_frame_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[40]_i_1_n_0 ,\pause_frame_good_reg[40]_i_1_n_1 ,\pause_frame_good_reg[40]_i_1_n_2 ,\pause_frame_good_reg[40]_i_1_n_3 ,\pause_frame_good_reg[40]_i_1_n_4 ,\pause_frame_good_reg[40]_i_1_n_5 ,\pause_frame_good_reg[40]_i_1_n_6 ,\pause_frame_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[40]_i_1_n_8 ,\pause_frame_good_reg[40]_i_1_n_9 ,\pause_frame_good_reg[40]_i_1_n_10 ,\pause_frame_good_reg[40]_i_1_n_11 ,\pause_frame_good_reg[40]_i_1_n_12 ,\pause_frame_good_reg[40]_i_1_n_13 ,\pause_frame_good_reg[40]_i_1_n_14 ,\pause_frame_good_reg[40]_i_1_n_15 }),
        .S(pause_frame_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_14 ),
        .Q(pause_frame_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_13 ),
        .Q(pause_frame_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_12 ),
        .Q(pause_frame_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_11 ),
        .Q(pause_frame_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_10 ),
        .Q(pause_frame_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_9 ),
        .Q(pause_frame_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[40]_i_1_n_8 ),
        .Q(pause_frame_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_15 ),
        .Q(pause_frame_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[48]_i_1 
       (.CI(\pause_frame_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[48]_i_1_n_0 ,\pause_frame_good_reg[48]_i_1_n_1 ,\pause_frame_good_reg[48]_i_1_n_2 ,\pause_frame_good_reg[48]_i_1_n_3 ,\pause_frame_good_reg[48]_i_1_n_4 ,\pause_frame_good_reg[48]_i_1_n_5 ,\pause_frame_good_reg[48]_i_1_n_6 ,\pause_frame_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[48]_i_1_n_8 ,\pause_frame_good_reg[48]_i_1_n_9 ,\pause_frame_good_reg[48]_i_1_n_10 ,\pause_frame_good_reg[48]_i_1_n_11 ,\pause_frame_good_reg[48]_i_1_n_12 ,\pause_frame_good_reg[48]_i_1_n_13 ,\pause_frame_good_reg[48]_i_1_n_14 ,\pause_frame_good_reg[48]_i_1_n_15 }),
        .S(pause_frame_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_14 ),
        .Q(pause_frame_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_11 ),
        .Q(pause_frame_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_13 ),
        .Q(pause_frame_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_12 ),
        .Q(pause_frame_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_11 ),
        .Q(pause_frame_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_10 ),
        .Q(pause_frame_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_9 ),
        .Q(pause_frame_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[48]_i_1_n_8 ),
        .Q(pause_frame_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_15 ),
        .Q(pause_frame_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[56]_i_1 
       (.CI(\pause_frame_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_pause_frame_good_reg[56]_i_1_CO_UNCONNECTED [7],\pause_frame_good_reg[56]_i_1_n_1 ,\pause_frame_good_reg[56]_i_1_n_2 ,\pause_frame_good_reg[56]_i_1_n_3 ,\pause_frame_good_reg[56]_i_1_n_4 ,\pause_frame_good_reg[56]_i_1_n_5 ,\pause_frame_good_reg[56]_i_1_n_6 ,\pause_frame_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[56]_i_1_n_8 ,\pause_frame_good_reg[56]_i_1_n_9 ,\pause_frame_good_reg[56]_i_1_n_10 ,\pause_frame_good_reg[56]_i_1_n_11 ,\pause_frame_good_reg[56]_i_1_n_12 ,\pause_frame_good_reg[56]_i_1_n_13 ,\pause_frame_good_reg[56]_i_1_n_14 ,\pause_frame_good_reg[56]_i_1_n_15 }),
        .S(pause_frame_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_14 ),
        .Q(pause_frame_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_13 ),
        .Q(pause_frame_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_12 ),
        .Q(pause_frame_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_10 ),
        .Q(pause_frame_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_11 ),
        .Q(pause_frame_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_10 ),
        .Q(pause_frame_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_9 ),
        .Q(pause_frame_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[56]_i_1_n_8 ),
        .Q(pause_frame_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_9 ),
        .Q(pause_frame_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[0]_i_1_n_8 ),
        .Q(pause_frame_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_15 ),
        .Q(pause_frame_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_good_reg[8]_i_1 
       (.CI(\pause_frame_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_good_reg[8]_i_1_n_0 ,\pause_frame_good_reg[8]_i_1_n_1 ,\pause_frame_good_reg[8]_i_1_n_2 ,\pause_frame_good_reg[8]_i_1_n_3 ,\pause_frame_good_reg[8]_i_1_n_4 ,\pause_frame_good_reg[8]_i_1_n_5 ,\pause_frame_good_reg[8]_i_1_n_6 ,\pause_frame_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_good_reg[8]_i_1_n_8 ,\pause_frame_good_reg[8]_i_1_n_9 ,\pause_frame_good_reg[8]_i_1_n_10 ,\pause_frame_good_reg[8]_i_1_n_11 ,\pause_frame_good_reg[8]_i_1_n_12 ,\pause_frame_good_reg[8]_i_1_n_13 ,\pause_frame_good_reg[8]_i_1_n_14 ,\pause_frame_good_reg[8]_i_1_n_15 }),
        .S(pause_frame_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_good_reg[8]_i_1_n_14 ),
        .Q(pause_frame_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \pause_frame_transed[0]_i_2 
       (.I0(pause_frame_transed_reg[0]),
        .O(\pause_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[0]_i_1_n_0 ,\pause_frame_transed_reg[0]_i_1_n_1 ,\pause_frame_transed_reg[0]_i_1_n_2 ,\pause_frame_transed_reg[0]_i_1_n_3 ,\pause_frame_transed_reg[0]_i_1_n_4 ,\pause_frame_transed_reg[0]_i_1_n_5 ,\pause_frame_transed_reg[0]_i_1_n_6 ,\pause_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\pause_frame_transed_reg[0]_i_1_n_8 ,\pause_frame_transed_reg[0]_i_1_n_9 ,\pause_frame_transed_reg[0]_i_1_n_10 ,\pause_frame_transed_reg[0]_i_1_n_11 ,\pause_frame_transed_reg[0]_i_1_n_12 ,\pause_frame_transed_reg[0]_i_1_n_13 ,\pause_frame_transed_reg[0]_i_1_n_14 ,\pause_frame_transed_reg[0]_i_1_n_15 }),
        .S({pause_frame_transed_reg[7:1],\pause_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[16]_i_1 
       (.CI(\pause_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[16]_i_1_n_0 ,\pause_frame_transed_reg[16]_i_1_n_1 ,\pause_frame_transed_reg[16]_i_1_n_2 ,\pause_frame_transed_reg[16]_i_1_n_3 ,\pause_frame_transed_reg[16]_i_1_n_4 ,\pause_frame_transed_reg[16]_i_1_n_5 ,\pause_frame_transed_reg[16]_i_1_n_6 ,\pause_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[16]_i_1_n_8 ,\pause_frame_transed_reg[16]_i_1_n_9 ,\pause_frame_transed_reg[16]_i_1_n_10 ,\pause_frame_transed_reg[16]_i_1_n_11 ,\pause_frame_transed_reg[16]_i_1_n_12 ,\pause_frame_transed_reg[16]_i_1_n_13 ,\pause_frame_transed_reg[16]_i_1_n_14 ,\pause_frame_transed_reg[16]_i_1_n_15 }),
        .S(pause_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[16]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[24]_i_1 
       (.CI(\pause_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[24]_i_1_n_0 ,\pause_frame_transed_reg[24]_i_1_n_1 ,\pause_frame_transed_reg[24]_i_1_n_2 ,\pause_frame_transed_reg[24]_i_1_n_3 ,\pause_frame_transed_reg[24]_i_1_n_4 ,\pause_frame_transed_reg[24]_i_1_n_5 ,\pause_frame_transed_reg[24]_i_1_n_6 ,\pause_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[24]_i_1_n_8 ,\pause_frame_transed_reg[24]_i_1_n_9 ,\pause_frame_transed_reg[24]_i_1_n_10 ,\pause_frame_transed_reg[24]_i_1_n_11 ,\pause_frame_transed_reg[24]_i_1_n_12 ,\pause_frame_transed_reg[24]_i_1_n_13 ,\pause_frame_transed_reg[24]_i_1_n_14 ,\pause_frame_transed_reg[24]_i_1_n_15 }),
        .S(pause_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[24]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[32]_i_1 
       (.CI(\pause_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[32]_i_1_n_0 ,\pause_frame_transed_reg[32]_i_1_n_1 ,\pause_frame_transed_reg[32]_i_1_n_2 ,\pause_frame_transed_reg[32]_i_1_n_3 ,\pause_frame_transed_reg[32]_i_1_n_4 ,\pause_frame_transed_reg[32]_i_1_n_5 ,\pause_frame_transed_reg[32]_i_1_n_6 ,\pause_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[32]_i_1_n_8 ,\pause_frame_transed_reg[32]_i_1_n_9 ,\pause_frame_transed_reg[32]_i_1_n_10 ,\pause_frame_transed_reg[32]_i_1_n_11 ,\pause_frame_transed_reg[32]_i_1_n_12 ,\pause_frame_transed_reg[32]_i_1_n_13 ,\pause_frame_transed_reg[32]_i_1_n_14 ,\pause_frame_transed_reg[32]_i_1_n_15 }),
        .S(pause_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[32]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[40]_i_1 
       (.CI(\pause_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[40]_i_1_n_0 ,\pause_frame_transed_reg[40]_i_1_n_1 ,\pause_frame_transed_reg[40]_i_1_n_2 ,\pause_frame_transed_reg[40]_i_1_n_3 ,\pause_frame_transed_reg[40]_i_1_n_4 ,\pause_frame_transed_reg[40]_i_1_n_5 ,\pause_frame_transed_reg[40]_i_1_n_6 ,\pause_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[40]_i_1_n_8 ,\pause_frame_transed_reg[40]_i_1_n_9 ,\pause_frame_transed_reg[40]_i_1_n_10 ,\pause_frame_transed_reg[40]_i_1_n_11 ,\pause_frame_transed_reg[40]_i_1_n_12 ,\pause_frame_transed_reg[40]_i_1_n_13 ,\pause_frame_transed_reg[40]_i_1_n_14 ,\pause_frame_transed_reg[40]_i_1_n_15 }),
        .S(pause_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[40]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[48]_i_1 
       (.CI(\pause_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[48]_i_1_n_0 ,\pause_frame_transed_reg[48]_i_1_n_1 ,\pause_frame_transed_reg[48]_i_1_n_2 ,\pause_frame_transed_reg[48]_i_1_n_3 ,\pause_frame_transed_reg[48]_i_1_n_4 ,\pause_frame_transed_reg[48]_i_1_n_5 ,\pause_frame_transed_reg[48]_i_1_n_6 ,\pause_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[48]_i_1_n_8 ,\pause_frame_transed_reg[48]_i_1_n_9 ,\pause_frame_transed_reg[48]_i_1_n_10 ,\pause_frame_transed_reg[48]_i_1_n_11 ,\pause_frame_transed_reg[48]_i_1_n_12 ,\pause_frame_transed_reg[48]_i_1_n_13 ,\pause_frame_transed_reg[48]_i_1_n_14 ,\pause_frame_transed_reg[48]_i_1_n_15 }),
        .S(pause_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[48]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[56]_i_1 
       (.CI(\pause_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_pause_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\pause_frame_transed_reg[56]_i_1_n_1 ,\pause_frame_transed_reg[56]_i_1_n_2 ,\pause_frame_transed_reg[56]_i_1_n_3 ,\pause_frame_transed_reg[56]_i_1_n_4 ,\pause_frame_transed_reg[56]_i_1_n_5 ,\pause_frame_transed_reg[56]_i_1_n_6 ,\pause_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[56]_i_1_n_8 ,\pause_frame_transed_reg[56]_i_1_n_9 ,\pause_frame_transed_reg[56]_i_1_n_10 ,\pause_frame_transed_reg[56]_i_1_n_11 ,\pause_frame_transed_reg[56]_i_1_n_12 ,\pause_frame_transed_reg[56]_i_1_n_13 ,\pause_frame_transed_reg[56]_i_1_n_14 ,\pause_frame_transed_reg[56]_i_1_n_15 }),
        .S(pause_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_13 ),
        .Q(pause_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_12 ),
        .Q(pause_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_11 ),
        .Q(pause_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_10 ),
        .Q(pause_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[56]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_9 ),
        .Q(pause_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[0]_i_1_n_8 ),
        .Q(pause_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_15 ),
        .Q(pause_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \pause_frame_transed_reg[8]_i_1 
       (.CI(\pause_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\pause_frame_transed_reg[8]_i_1_n_0 ,\pause_frame_transed_reg[8]_i_1_n_1 ,\pause_frame_transed_reg[8]_i_1_n_2 ,\pause_frame_transed_reg[8]_i_1_n_3 ,\pause_frame_transed_reg[8]_i_1_n_4 ,\pause_frame_transed_reg[8]_i_1_n_5 ,\pause_frame_transed_reg[8]_i_1_n_6 ,\pause_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\pause_frame_transed_reg[8]_i_1_n_8 ,\pause_frame_transed_reg[8]_i_1_n_9 ,\pause_frame_transed_reg[8]_i_1_n_10 ,\pause_frame_transed_reg[8]_i_1_n_11 ,\pause_frame_transed_reg[8]_i_1_n_12 ,\pause_frame_transed_reg[8]_i_1_n_13 ,\pause_frame_transed_reg[8]_i_1_n_14 ,\pause_frame_transed_reg[8]_i_1_n_15 }),
        .S(pause_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \pause_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[13]),
        .CLR(rst_i),
        .D(\pause_frame_transed_reg[8]_i_1_n_14 ),
        .Q(pause_frame_transed_reg[9]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h8)) 
    read_done_i_1
       (.I0(\state_reg_n_0_[1] ),
        .I1(data_sel),
        .O(read_done_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    read_done_reg
       (.C(clk_i),
        .CE(read_done),
        .CLR(rst_i),
        .D(read_done_i_1_n_0),
        .Q(read_done_reg_n_0));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \recv_config0[31]_i_1 
       (.I0(\recv_config0_reg[0]_0 ),
        .I1(out[9]),
        .I2(\stat_rd_data_reg[63]_1 ),
        .I3(\recv_config0[31]_i_2_n_0 ),
        .I4(\recv_config0[31]_i_3_n_0 ),
        .I5(out[7]),
        .O(\recv_config0[31]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \recv_config0[31]_i_2 
       (.I0(out[6]),
        .I1(out[8]),
        .I2(out[4]),
        .I3(out[5]),
        .O(\recv_config0[31]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \recv_config0[31]_i_3 
       (.I0(out[2]),
        .I1(out[3]),
        .I2(out[0]),
        .I3(out[1]),
        .O(\recv_config0[31]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[0] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[0]),
        .Q(cfgRxRegData[0]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[10] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[10]),
        .Q(cfgRxRegData[10]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[11] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[11]),
        .Q(cfgRxRegData[11]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[12] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[12]),
        .Q(cfgRxRegData[12]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[13] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[13]),
        .Q(cfgRxRegData[13]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[14] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[14]),
        .Q(cfgRxRegData[14]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[15] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[15]),
        .Q(cfgRxRegData[15]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[16] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[16]),
        .Q(cfgRxRegData[16]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[17] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[17]),
        .Q(cfgRxRegData[17]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[18] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[18]),
        .Q(cfgRxRegData[18]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[19] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[19]),
        .Q(cfgRxRegData[19]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[1] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[1]),
        .Q(cfgRxRegData[1]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[20] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[20]),
        .Q(cfgRxRegData[20]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[21] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[21]),
        .Q(cfgRxRegData[21]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[22] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[22]),
        .Q(cfgRxRegData[22]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[23] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[23]),
        .Q(cfgRxRegData[23]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[24] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[24]),
        .Q(cfgRxRegData[24]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[25] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[25]),
        .Q(cfgRxRegData[25]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[26] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[26]),
        .Q(cfgRxRegData[26]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[27] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[27]),
        .Q(cfgRxRegData[27]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[28] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[28]),
        .Q(cfgRxRegData[28]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[29] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[29]),
        .Q(cfgRxRegData[29]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[2] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[2]),
        .Q(cfgRxRegData[2]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[30] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[30]),
        .Q(cfgRxRegData[30]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[31] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[31]),
        .Q(cfgRxRegData[31]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[3] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[3]),
        .Q(cfgRxRegData[3]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[4] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[4]),
        .Q(cfgRxRegData[4]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[5] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[5]),
        .Q(cfgRxRegData[5]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[6] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[6]),
        .Q(cfgRxRegData[6]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[7] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[7]),
        .Q(cfgRxRegData[7]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[8] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[8]),
        .Q(cfgRxRegData[8]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config0_reg[9] 
       (.C(clk_i),
        .CE(\recv_config0[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[9]),
        .Q(cfgRxRegData[9]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \recv_config1[31]_i_1 
       (.I0(recv_config01__0),
        .I1(\recv_config1[31]_i_3_n_0 ),
        .I2(out[7]),
        .I3(out[8]),
        .I4(\recv_config1[31]_i_4_n_0 ),
        .I5(out[6]),
        .O(\recv_config1[31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \recv_config1[31]_i_2 
       (.I0(\stat_rd_data_reg[63]_1 ),
        .I1(out[9]),
        .I2(\recv_config0_reg[0]_0 ),
        .O(recv_config01__0));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \recv_config1[31]_i_3 
       (.I0(out[0]),
        .I1(out[5]),
        .O(\recv_config1[31]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \recv_config1[31]_i_4 
       (.I0(out[3]),
        .I1(out[4]),
        .I2(out[1]),
        .I3(out[2]),
        .O(\recv_config1[31]_i_4_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[0] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[0]),
        .Q(cfgRxRegData[32]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[10] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[10]),
        .Q(cfgRxRegData[42]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[11] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[11]),
        .Q(cfgRxRegData[43]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[12] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[12]),
        .Q(cfgRxRegData[44]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[13] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[13]),
        .Q(cfgRxRegData[45]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[14] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[14]),
        .Q(cfgRxRegData[46]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[15] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[15]),
        .Q(cfgRxRegData[47]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[16] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[16]),
        .Q(\recv_config1_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[17] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[17]),
        .Q(\recv_config1_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[18] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[18]),
        .Q(\recv_config1_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[19] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[19]),
        .Q(\recv_config1_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[1] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[1]),
        .Q(cfgRxRegData[33]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[20] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[20]),
        .Q(\recv_config1_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[21] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[21]),
        .Q(\recv_config1_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[22] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[22]),
        .Q(\recv_config1_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[23] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[23]),
        .Q(\recv_config1_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[24] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[24]),
        .Q(\recv_config1_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[25] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[25]),
        .Q(\recv_config1_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[26] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[26]),
        .Q(\recv_config1_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[27] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[27]),
        .Q(cfgRxRegData[48]));
  FDPE #(
    .INIT(1'b1)) 
    \recv_config1_reg[28] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .D(mgmt_wr_data[28]),
        .PRE(rst_i),
        .Q(cfgRxRegData[49]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[29] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[29]),
        .Q(cfgRxRegData[50]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[2] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[2]),
        .Q(cfgRxRegData[34]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[30] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[30]),
        .Q(cfgRxRegData[51]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[31] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[31]),
        .Q(cfgRxRegData[52]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[3] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[3]),
        .Q(cfgRxRegData[35]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[4] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[4]),
        .Q(cfgRxRegData[36]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[5] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[5]),
        .Q(cfgRxRegData[37]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[6] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[6]),
        .Q(cfgRxRegData[38]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[7] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[7]),
        .Q(cfgRxRegData[39]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[8] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[8]),
        .Q(cfgRxRegData[40]));
  FDCE #(
    .INIT(1'b0)) 
    \recv_config1_reg[9] 
       (.C(clk_i),
        .CE(\recv_config1[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[9]),
        .Q(cfgRxRegData[41]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \rs_config[31]_i_1 
       (.I0(\recv_config0_reg[0]_0 ),
        .I1(out[9]),
        .I2(\stat_rd_data_reg[63]_1 ),
        .I3(\rs_config[31]_i_2_n_0 ),
        .I4(\recv_config1[31]_i_4_n_0 ),
        .I5(out[8]),
        .O(\rs_config[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rs_config[31]_i_2 
       (.I0(out[0]),
        .I1(out[7]),
        .I2(out[5]),
        .I3(out[6]),
        .O(\rs_config[31]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[0] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[0]),
        .Q(\rs_config_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[10] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[10]),
        .Q(\rs_config_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[11] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[11]),
        .Q(\rs_config_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[12] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[12]),
        .Q(\rs_config_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[13] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[13]),
        .Q(\rs_config_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[14] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[14]),
        .Q(\rs_config_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[15] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[15]),
        .Q(\rs_config_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[16] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[16]),
        .Q(\rs_config_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[17] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[17]),
        .Q(\rs_config_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[18] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[18]),
        .Q(\rs_config_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[19] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[19]),
        .Q(\rs_config_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[1] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[1]),
        .Q(\rs_config_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[20] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[20]),
        .Q(\rs_config_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[21] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[21]),
        .Q(\rs_config_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[22] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[22]),
        .Q(\rs_config_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[23] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[23]),
        .Q(\rs_config_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[24] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[24]),
        .Q(\rs_config_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[25] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[25]),
        .Q(\rs_config_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[26] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[26]),
        .Q(\rs_config_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[27] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[27]),
        .Q(cfgTxRegData[9]));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[28] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[28]),
        .Q(\rs_config_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[29] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[29]),
        .Q(\rs_config_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[2] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[2]),
        .Q(\rs_config_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[30] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[30]),
        .Q(\rs_config_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[31] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[31]),
        .Q(\rs_config_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[3] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[3]),
        .Q(\rs_config_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[4] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[4]),
        .Q(\rs_config_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[5] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[5]),
        .Q(\rs_config_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[6] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[6]),
        .Q(\rs_config_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[7] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[7]),
        .Q(\rs_config_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[8] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[8]),
        .Q(\rs_config_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \rs_config_reg[9] 
       (.C(clk_i),
        .CE(\rs_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[9]),
        .Q(\rs_config_reg_n_0_[9] ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[0]_i_1 
       (.I0(\stat_rd_data[0]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[0]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_10 
       (.I0(tagged_frame_transed_reg[0]),
        .I1(frame_1024_max_transed_reg[0]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[0]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[0]),
        .O(\stat_rd_data[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_11 
       (.I0(multicast_received_good_reg[0]),
        .I1(broadcast_received_good_reg[0]),
        .I2(out[1]),
        .I3(fcs_error_reg[0]),
        .I4(out[0]),
        .I5(frame_received_good_reg[0]),
        .O(\stat_rd_data[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_12 
       (.I0(frame_256_511_good_reg[0]),
        .I1(frame_128_255_good_reg[0]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[0]),
        .I4(out[0]),
        .I5(frame_64_good_reg[0]),
        .O(\stat_rd_data[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_13 
       (.I0(lt_out_range_reg[0]),
        .I1(control_frame_good_reg[0]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[0]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[0]),
        .O(\stat_rd_data[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_14 
       (.I0(oversize_frame_good_reg[0]),
        .I1(unsupported_control_frame_reg[0]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[0]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[0]),
        .O(\stat_rd_data[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_2 
       (.I0(\stat_rd_data_reg[0]_i_4_n_0 ),
        .I1(\stat_rd_data[0]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[0]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[0]_i_7_n_0 ),
        .O(\stat_rd_data[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_3 
       (.I0(total_bytes_transed_reg[0]),
        .I1(total_bytes_recved_reg[0]),
        .I2(out[1]),
        .I3(fragment_frame_reg[0]),
        .I4(out[0]),
        .I5(undersize_frame_reg[0]),
        .O(\stat_rd_data[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[0]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[0]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[0]),
        .I5(pause_frame_transed_reg[0]),
        .O(\stat_rd_data[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_6 
       (.I0(frame_128_255_transed_reg[0]),
        .I1(frame_65_127_transed_reg[0]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[0]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[0]),
        .O(\stat_rd_data[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[0]_i_7 
       (.I0(underrun_error_reg[0]),
        .I1(multicast_frame_transed_reg[0]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[0]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[0]),
        .O(\stat_rd_data[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[10]_i_1 
       (.I0(\stat_rd_data[10]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[10]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_10 
       (.I0(tagged_frame_transed_reg[10]),
        .I1(frame_1024_max_transed_reg[10]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[10]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[10]),
        .O(\stat_rd_data[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_11 
       (.I0(multicast_received_good_reg[10]),
        .I1(broadcast_received_good_reg[10]),
        .I2(out[1]),
        .I3(fcs_error_reg[10]),
        .I4(out[0]),
        .I5(frame_received_good_reg[10]),
        .O(\stat_rd_data[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_12 
       (.I0(frame_256_511_good_reg[10]),
        .I1(frame_128_255_good_reg[10]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[10]),
        .I4(out[0]),
        .I5(frame_64_good_reg[10]),
        .O(\stat_rd_data[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_13 
       (.I0(lt_out_range_reg[10]),
        .I1(control_frame_good_reg[10]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[10]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[10]),
        .O(\stat_rd_data[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_14 
       (.I0(oversize_frame_good_reg[10]),
        .I1(unsupported_control_frame_reg[10]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[10]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[10]),
        .O(\stat_rd_data[10]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_2 
       (.I0(\stat_rd_data_reg[10]_i_4_n_0 ),
        .I1(\stat_rd_data[10]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[10]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[10]_i_7_n_0 ),
        .O(\stat_rd_data[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_3 
       (.I0(total_bytes_transed_reg[10]),
        .I1(total_bytes_recved_reg[10]),
        .I2(out[1]),
        .I3(fragment_frame_reg[10]),
        .I4(out[0]),
        .I5(undersize_frame_reg[10]),
        .O(\stat_rd_data[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[10]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[10]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[10]),
        .I5(pause_frame_transed_reg[10]),
        .O(\stat_rd_data[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_6 
       (.I0(frame_128_255_transed_reg[10]),
        .I1(frame_65_127_transed_reg[10]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[10]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[10]),
        .O(\stat_rd_data[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[10]_i_7 
       (.I0(underrun_error_reg[10]),
        .I1(multicast_frame_transed_reg[10]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[10]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[10]),
        .O(\stat_rd_data[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[11]_i_1 
       (.I0(\stat_rd_data[11]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[11]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_10 
       (.I0(tagged_frame_transed_reg[11]),
        .I1(frame_1024_max_transed_reg[11]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[11]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[11]),
        .O(\stat_rd_data[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_11 
       (.I0(multicast_received_good_reg[11]),
        .I1(broadcast_received_good_reg[11]),
        .I2(out[1]),
        .I3(fcs_error_reg[11]),
        .I4(out[0]),
        .I5(frame_received_good_reg[11]),
        .O(\stat_rd_data[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_12 
       (.I0(frame_256_511_good_reg[11]),
        .I1(frame_128_255_good_reg[11]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[11]),
        .I4(out[0]),
        .I5(frame_64_good_reg[11]),
        .O(\stat_rd_data[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_13 
       (.I0(lt_out_range_reg[11]),
        .I1(control_frame_good_reg[11]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[11]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[11]),
        .O(\stat_rd_data[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_14 
       (.I0(oversize_frame_good_reg[11]),
        .I1(unsupported_control_frame_reg[11]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[11]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[11]),
        .O(\stat_rd_data[11]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_2 
       (.I0(\stat_rd_data_reg[11]_i_4_n_0 ),
        .I1(\stat_rd_data[11]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[11]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[11]_i_7_n_0 ),
        .O(\stat_rd_data[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_3 
       (.I0(total_bytes_transed_reg[11]),
        .I1(total_bytes_recved_reg[11]),
        .I2(out[1]),
        .I3(fragment_frame_reg[11]),
        .I4(out[0]),
        .I5(undersize_frame_reg[11]),
        .O(\stat_rd_data[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[11]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[11]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[11]),
        .I5(pause_frame_transed_reg[11]),
        .O(\stat_rd_data[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_6 
       (.I0(frame_128_255_transed_reg[11]),
        .I1(frame_65_127_transed_reg[11]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[11]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[11]),
        .O(\stat_rd_data[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[11]_i_7 
       (.I0(underrun_error_reg[11]),
        .I1(multicast_frame_transed_reg[11]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[11]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[11]),
        .O(\stat_rd_data[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[12]_i_1 
       (.I0(\stat_rd_data[12]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[12]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_10 
       (.I0(tagged_frame_transed_reg[12]),
        .I1(frame_1024_max_transed_reg[12]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[12]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[12]),
        .O(\stat_rd_data[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_11 
       (.I0(multicast_received_good_reg[12]),
        .I1(broadcast_received_good_reg[12]),
        .I2(out[1]),
        .I3(fcs_error_reg[12]),
        .I4(out[0]),
        .I5(frame_received_good_reg[12]),
        .O(\stat_rd_data[12]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_12 
       (.I0(frame_256_511_good_reg[12]),
        .I1(frame_128_255_good_reg[12]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[12]),
        .I4(out[0]),
        .I5(frame_64_good_reg[12]),
        .O(\stat_rd_data[12]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_13 
       (.I0(lt_out_range_reg[12]),
        .I1(control_frame_good_reg[12]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[12]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[12]),
        .O(\stat_rd_data[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_14 
       (.I0(oversize_frame_good_reg[12]),
        .I1(unsupported_control_frame_reg[12]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[12]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[12]),
        .O(\stat_rd_data[12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_2 
       (.I0(\stat_rd_data_reg[12]_i_4_n_0 ),
        .I1(\stat_rd_data[12]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[12]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[12]_i_7_n_0 ),
        .O(\stat_rd_data[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_3 
       (.I0(total_bytes_transed_reg[12]),
        .I1(total_bytes_recved_reg[12]),
        .I2(out[1]),
        .I3(fragment_frame_reg[12]),
        .I4(out[0]),
        .I5(undersize_frame_reg[12]),
        .O(\stat_rd_data[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[12]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[12]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[12]),
        .I5(pause_frame_transed_reg[12]),
        .O(\stat_rd_data[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_6 
       (.I0(frame_128_255_transed_reg[12]),
        .I1(frame_65_127_transed_reg[12]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[12]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[12]),
        .O(\stat_rd_data[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[12]_i_7 
       (.I0(underrun_error_reg[12]),
        .I1(multicast_frame_transed_reg[12]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[12]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[12]),
        .O(\stat_rd_data[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[13]_i_1 
       (.I0(\stat_rd_data[13]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[13]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_10 
       (.I0(tagged_frame_transed_reg[13]),
        .I1(frame_1024_max_transed_reg[13]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[13]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[13]),
        .O(\stat_rd_data[13]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_11 
       (.I0(multicast_received_good_reg[13]),
        .I1(broadcast_received_good_reg[13]),
        .I2(out[1]),
        .I3(fcs_error_reg[13]),
        .I4(out[0]),
        .I5(frame_received_good_reg[13]),
        .O(\stat_rd_data[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_12 
       (.I0(frame_256_511_good_reg[13]),
        .I1(frame_128_255_good_reg[13]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[13]),
        .I4(out[0]),
        .I5(frame_64_good_reg[13]),
        .O(\stat_rd_data[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_13 
       (.I0(lt_out_range_reg[13]),
        .I1(control_frame_good_reg[13]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[13]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[13]),
        .O(\stat_rd_data[13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_14 
       (.I0(oversize_frame_good_reg[13]),
        .I1(unsupported_control_frame_reg[13]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[13]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[13]),
        .O(\stat_rd_data[13]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_2 
       (.I0(\stat_rd_data_reg[13]_i_4_n_0 ),
        .I1(\stat_rd_data[13]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[13]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[13]_i_7_n_0 ),
        .O(\stat_rd_data[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_3 
       (.I0(total_bytes_transed_reg[13]),
        .I1(total_bytes_recved_reg[13]),
        .I2(out[1]),
        .I3(fragment_frame_reg[13]),
        .I4(out[0]),
        .I5(undersize_frame_reg[13]),
        .O(\stat_rd_data[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[13]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[13]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[13]),
        .I5(pause_frame_transed_reg[13]),
        .O(\stat_rd_data[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_6 
       (.I0(frame_128_255_transed_reg[13]),
        .I1(frame_65_127_transed_reg[13]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[13]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[13]),
        .O(\stat_rd_data[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[13]_i_7 
       (.I0(underrun_error_reg[13]),
        .I1(multicast_frame_transed_reg[13]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[13]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[13]),
        .O(\stat_rd_data[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[14]_i_1 
       (.I0(\stat_rd_data[14]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[14]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_10 
       (.I0(tagged_frame_transed_reg[14]),
        .I1(frame_1024_max_transed_reg[14]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[14]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[14]),
        .O(\stat_rd_data[14]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_11 
       (.I0(multicast_received_good_reg[14]),
        .I1(broadcast_received_good_reg[14]),
        .I2(out[1]),
        .I3(fcs_error_reg[14]),
        .I4(out[0]),
        .I5(frame_received_good_reg[14]),
        .O(\stat_rd_data[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_12 
       (.I0(frame_256_511_good_reg[14]),
        .I1(frame_128_255_good_reg[14]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[14]),
        .I4(out[0]),
        .I5(frame_64_good_reg[14]),
        .O(\stat_rd_data[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_13 
       (.I0(lt_out_range_reg[14]),
        .I1(control_frame_good_reg[14]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[14]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[14]),
        .O(\stat_rd_data[14]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_14 
       (.I0(oversize_frame_good_reg[14]),
        .I1(unsupported_control_frame_reg[14]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[14]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[14]),
        .O(\stat_rd_data[14]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_2 
       (.I0(\stat_rd_data_reg[14]_i_4_n_0 ),
        .I1(\stat_rd_data[14]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[14]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[14]_i_7_n_0 ),
        .O(\stat_rd_data[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_3 
       (.I0(total_bytes_transed_reg[14]),
        .I1(total_bytes_recved_reg[14]),
        .I2(out[1]),
        .I3(fragment_frame_reg[14]),
        .I4(out[0]),
        .I5(undersize_frame_reg[14]),
        .O(\stat_rd_data[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[14]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[14]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[14]),
        .I5(pause_frame_transed_reg[14]),
        .O(\stat_rd_data[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_6 
       (.I0(frame_128_255_transed_reg[14]),
        .I1(frame_65_127_transed_reg[14]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[14]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[14]),
        .O(\stat_rd_data[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[14]_i_7 
       (.I0(underrun_error_reg[14]),
        .I1(multicast_frame_transed_reg[14]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[14]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[14]),
        .O(\stat_rd_data[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[15]_i_1 
       (.I0(\stat_rd_data[15]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[15]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_10 
       (.I0(tagged_frame_transed_reg[15]),
        .I1(frame_1024_max_transed_reg[15]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[15]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[15]),
        .O(\stat_rd_data[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_11 
       (.I0(multicast_received_good_reg[15]),
        .I1(broadcast_received_good_reg[15]),
        .I2(out[1]),
        .I3(fcs_error_reg[15]),
        .I4(out[0]),
        .I5(frame_received_good_reg[15]),
        .O(\stat_rd_data[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_12 
       (.I0(frame_256_511_good_reg[15]),
        .I1(frame_128_255_good_reg[15]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[15]),
        .I4(out[0]),
        .I5(frame_64_good_reg[15]),
        .O(\stat_rd_data[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_13 
       (.I0(lt_out_range_reg[15]),
        .I1(control_frame_good_reg[15]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[15]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[15]),
        .O(\stat_rd_data[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_14 
       (.I0(oversize_frame_good_reg[15]),
        .I1(unsupported_control_frame_reg[15]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[15]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[15]),
        .O(\stat_rd_data[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_2 
       (.I0(\stat_rd_data_reg[15]_i_4_n_0 ),
        .I1(\stat_rd_data[15]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[15]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[15]_i_7_n_0 ),
        .O(\stat_rd_data[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_3 
       (.I0(total_bytes_transed_reg[15]),
        .I1(total_bytes_recved_reg[15]),
        .I2(out[1]),
        .I3(fragment_frame_reg[15]),
        .I4(out[0]),
        .I5(undersize_frame_reg[15]),
        .O(\stat_rd_data[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[15]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[15]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[15]),
        .I5(pause_frame_transed_reg[15]),
        .O(\stat_rd_data[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_6 
       (.I0(frame_128_255_transed_reg[15]),
        .I1(frame_65_127_transed_reg[15]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[15]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[15]),
        .O(\stat_rd_data[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[15]_i_7 
       (.I0(underrun_error_reg[15]),
        .I1(multicast_frame_transed_reg[15]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[15]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[15]),
        .O(\stat_rd_data[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[16]_i_1 
       (.I0(\stat_rd_data[16]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[16]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_10 
       (.I0(tagged_frame_transed_reg[16]),
        .I1(frame_1024_max_transed_reg[16]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[16]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[16]),
        .O(\stat_rd_data[16]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_11 
       (.I0(multicast_received_good_reg[16]),
        .I1(broadcast_received_good_reg[16]),
        .I2(out[1]),
        .I3(fcs_error_reg[16]),
        .I4(out[0]),
        .I5(frame_received_good_reg[16]),
        .O(\stat_rd_data[16]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_12 
       (.I0(frame_256_511_good_reg[16]),
        .I1(frame_128_255_good_reg[16]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[16]),
        .I4(out[0]),
        .I5(frame_64_good_reg[16]),
        .O(\stat_rd_data[16]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_13 
       (.I0(lt_out_range_reg[16]),
        .I1(control_frame_good_reg[16]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[16]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[16]),
        .O(\stat_rd_data[16]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_14 
       (.I0(oversize_frame_good_reg[16]),
        .I1(unsupported_control_frame_reg[16]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[16]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[16]),
        .O(\stat_rd_data[16]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_2 
       (.I0(\stat_rd_data_reg[16]_i_4_n_0 ),
        .I1(\stat_rd_data[16]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[16]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[16]_i_7_n_0 ),
        .O(\stat_rd_data[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_3 
       (.I0(total_bytes_transed_reg[16]),
        .I1(total_bytes_recved_reg[16]),
        .I2(out[1]),
        .I3(fragment_frame_reg[16]),
        .I4(out[0]),
        .I5(undersize_frame_reg[16]),
        .O(\stat_rd_data[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[16]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[16]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[16]),
        .I5(pause_frame_transed_reg[16]),
        .O(\stat_rd_data[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_6 
       (.I0(frame_128_255_transed_reg[16]),
        .I1(frame_65_127_transed_reg[16]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[16]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[16]),
        .O(\stat_rd_data[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[16]_i_7 
       (.I0(underrun_error_reg[16]),
        .I1(multicast_frame_transed_reg[16]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[16]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[16]),
        .O(\stat_rd_data[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[17]_i_1 
       (.I0(\stat_rd_data[17]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[17]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[17]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_10 
       (.I0(tagged_frame_transed_reg[17]),
        .I1(frame_1024_max_transed_reg[17]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[17]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[17]),
        .O(\stat_rd_data[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_11 
       (.I0(multicast_received_good_reg[17]),
        .I1(broadcast_received_good_reg[17]),
        .I2(out[1]),
        .I3(fcs_error_reg[17]),
        .I4(out[0]),
        .I5(frame_received_good_reg[17]),
        .O(\stat_rd_data[17]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_12 
       (.I0(frame_256_511_good_reg[17]),
        .I1(frame_128_255_good_reg[17]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[17]),
        .I4(out[0]),
        .I5(frame_64_good_reg[17]),
        .O(\stat_rd_data[17]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_13 
       (.I0(lt_out_range_reg[17]),
        .I1(control_frame_good_reg[17]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[17]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[17]),
        .O(\stat_rd_data[17]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_14 
       (.I0(oversize_frame_good_reg[17]),
        .I1(unsupported_control_frame_reg[17]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[17]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[17]),
        .O(\stat_rd_data[17]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_2 
       (.I0(\stat_rd_data_reg[17]_i_4_n_0 ),
        .I1(\stat_rd_data[17]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[17]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[17]_i_7_n_0 ),
        .O(\stat_rd_data[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_3 
       (.I0(total_bytes_transed_reg[17]),
        .I1(total_bytes_recved_reg[17]),
        .I2(out[1]),
        .I3(fragment_frame_reg[17]),
        .I4(out[0]),
        .I5(undersize_frame_reg[17]),
        .O(\stat_rd_data[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[17]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[17]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[17]),
        .I5(pause_frame_transed_reg[17]),
        .O(\stat_rd_data[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_6 
       (.I0(frame_128_255_transed_reg[17]),
        .I1(frame_65_127_transed_reg[17]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[17]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[17]),
        .O(\stat_rd_data[17]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[17]_i_7 
       (.I0(underrun_error_reg[17]),
        .I1(multicast_frame_transed_reg[17]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[17]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[17]),
        .O(\stat_rd_data[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[18]_i_1 
       (.I0(\stat_rd_data[18]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[18]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_10 
       (.I0(tagged_frame_transed_reg[18]),
        .I1(frame_1024_max_transed_reg[18]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[18]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[18]),
        .O(\stat_rd_data[18]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_11 
       (.I0(multicast_received_good_reg[18]),
        .I1(broadcast_received_good_reg[18]),
        .I2(out[1]),
        .I3(fcs_error_reg[18]),
        .I4(out[0]),
        .I5(frame_received_good_reg[18]),
        .O(\stat_rd_data[18]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_12 
       (.I0(frame_256_511_good_reg[18]),
        .I1(frame_128_255_good_reg[18]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[18]),
        .I4(out[0]),
        .I5(frame_64_good_reg[18]),
        .O(\stat_rd_data[18]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_13 
       (.I0(lt_out_range_reg[18]),
        .I1(control_frame_good_reg[18]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[18]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[18]),
        .O(\stat_rd_data[18]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_14 
       (.I0(oversize_frame_good_reg[18]),
        .I1(unsupported_control_frame_reg[18]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[18]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[18]),
        .O(\stat_rd_data[18]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_2 
       (.I0(\stat_rd_data_reg[18]_i_4_n_0 ),
        .I1(\stat_rd_data[18]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[18]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[18]_i_7_n_0 ),
        .O(\stat_rd_data[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_3 
       (.I0(total_bytes_transed_reg[18]),
        .I1(total_bytes_recved_reg[18]),
        .I2(out[1]),
        .I3(fragment_frame_reg[18]),
        .I4(out[0]),
        .I5(undersize_frame_reg[18]),
        .O(\stat_rd_data[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[18]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[18]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[18]),
        .I5(pause_frame_transed_reg[18]),
        .O(\stat_rd_data[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_6 
       (.I0(frame_128_255_transed_reg[18]),
        .I1(frame_65_127_transed_reg[18]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[18]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[18]),
        .O(\stat_rd_data[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[18]_i_7 
       (.I0(underrun_error_reg[18]),
        .I1(multicast_frame_transed_reg[18]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[18]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[18]),
        .O(\stat_rd_data[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[19]_i_1 
       (.I0(\stat_rd_data[19]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[19]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_10 
       (.I0(tagged_frame_transed_reg[19]),
        .I1(frame_1024_max_transed_reg[19]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[19]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[19]),
        .O(\stat_rd_data[19]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_11 
       (.I0(multicast_received_good_reg[19]),
        .I1(broadcast_received_good_reg[19]),
        .I2(out[1]),
        .I3(fcs_error_reg[19]),
        .I4(out[0]),
        .I5(frame_received_good_reg[19]),
        .O(\stat_rd_data[19]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_12 
       (.I0(frame_256_511_good_reg[19]),
        .I1(frame_128_255_good_reg[19]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[19]),
        .I4(out[0]),
        .I5(frame_64_good_reg[19]),
        .O(\stat_rd_data[19]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_13 
       (.I0(lt_out_range_reg[19]),
        .I1(control_frame_good_reg[19]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[19]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[19]),
        .O(\stat_rd_data[19]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_14 
       (.I0(oversize_frame_good_reg[19]),
        .I1(unsupported_control_frame_reg[19]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[19]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[19]),
        .O(\stat_rd_data[19]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_2 
       (.I0(\stat_rd_data_reg[19]_i_4_n_0 ),
        .I1(\stat_rd_data[19]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[19]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[19]_i_7_n_0 ),
        .O(\stat_rd_data[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_3 
       (.I0(total_bytes_transed_reg[19]),
        .I1(total_bytes_recved_reg[19]),
        .I2(out[1]),
        .I3(fragment_frame_reg[19]),
        .I4(out[0]),
        .I5(undersize_frame_reg[19]),
        .O(\stat_rd_data[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[19]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[19]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[19]),
        .I5(pause_frame_transed_reg[19]),
        .O(\stat_rd_data[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_6 
       (.I0(frame_128_255_transed_reg[19]),
        .I1(frame_65_127_transed_reg[19]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[19]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[19]),
        .O(\stat_rd_data[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[19]_i_7 
       (.I0(underrun_error_reg[19]),
        .I1(multicast_frame_transed_reg[19]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[19]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[19]),
        .O(\stat_rd_data[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[1]_i_1 
       (.I0(\stat_rd_data[1]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[1]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_10 
       (.I0(tagged_frame_transed_reg[1]),
        .I1(frame_1024_max_transed_reg[1]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[1]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[1]),
        .O(\stat_rd_data[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_11 
       (.I0(multicast_received_good_reg[1]),
        .I1(broadcast_received_good_reg[1]),
        .I2(out[1]),
        .I3(fcs_error_reg[1]),
        .I4(out[0]),
        .I5(frame_received_good_reg[1]),
        .O(\stat_rd_data[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_12 
       (.I0(frame_256_511_good_reg[1]),
        .I1(frame_128_255_good_reg[1]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[1]),
        .I4(out[0]),
        .I5(frame_64_good_reg[1]),
        .O(\stat_rd_data[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_13 
       (.I0(lt_out_range_reg[1]),
        .I1(control_frame_good_reg[1]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[1]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[1]),
        .O(\stat_rd_data[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_14 
       (.I0(oversize_frame_good_reg[1]),
        .I1(unsupported_control_frame_reg[1]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[1]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[1]),
        .O(\stat_rd_data[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_2 
       (.I0(\stat_rd_data_reg[1]_i_4_n_0 ),
        .I1(\stat_rd_data[1]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[1]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[1]_i_7_n_0 ),
        .O(\stat_rd_data[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_3 
       (.I0(total_bytes_transed_reg[1]),
        .I1(total_bytes_recved_reg[1]),
        .I2(out[1]),
        .I3(fragment_frame_reg[1]),
        .I4(out[0]),
        .I5(undersize_frame_reg[1]),
        .O(\stat_rd_data[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[1]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[1]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[1]),
        .I5(pause_frame_transed_reg[1]),
        .O(\stat_rd_data[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_6 
       (.I0(frame_128_255_transed_reg[1]),
        .I1(frame_65_127_transed_reg[1]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[1]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[1]),
        .O(\stat_rd_data[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[1]_i_7 
       (.I0(underrun_error_reg[1]),
        .I1(multicast_frame_transed_reg[1]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[1]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[1]),
        .O(\stat_rd_data[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[20]_i_1 
       (.I0(\stat_rd_data[20]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[20]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_10 
       (.I0(tagged_frame_transed_reg[20]),
        .I1(frame_1024_max_transed_reg[20]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[20]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[20]),
        .O(\stat_rd_data[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_11 
       (.I0(multicast_received_good_reg[20]),
        .I1(broadcast_received_good_reg[20]),
        .I2(out[1]),
        .I3(fcs_error_reg[20]),
        .I4(out[0]),
        .I5(frame_received_good_reg[20]),
        .O(\stat_rd_data[20]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_12 
       (.I0(frame_256_511_good_reg[20]),
        .I1(frame_128_255_good_reg[20]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[20]),
        .I4(out[0]),
        .I5(frame_64_good_reg[20]),
        .O(\stat_rd_data[20]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_13 
       (.I0(lt_out_range_reg[20]),
        .I1(control_frame_good_reg[20]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[20]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[20]),
        .O(\stat_rd_data[20]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_14 
       (.I0(oversize_frame_good_reg[20]),
        .I1(unsupported_control_frame_reg[20]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[20]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[20]),
        .O(\stat_rd_data[20]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_2 
       (.I0(\stat_rd_data_reg[20]_i_4_n_0 ),
        .I1(\stat_rd_data[20]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[20]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[20]_i_7_n_0 ),
        .O(\stat_rd_data[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_3 
       (.I0(total_bytes_transed_reg[20]),
        .I1(total_bytes_recved_reg[20]),
        .I2(out[1]),
        .I3(fragment_frame_reg[20]),
        .I4(out[0]),
        .I5(undersize_frame_reg[20]),
        .O(\stat_rd_data[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[20]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[20]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[20]),
        .I5(pause_frame_transed_reg[20]),
        .O(\stat_rd_data[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_6 
       (.I0(frame_128_255_transed_reg[20]),
        .I1(frame_65_127_transed_reg[20]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[20]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[20]),
        .O(\stat_rd_data[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[20]_i_7 
       (.I0(underrun_error_reg[20]),
        .I1(multicast_frame_transed_reg[20]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[20]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[20]),
        .O(\stat_rd_data[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[21]_i_1 
       (.I0(\stat_rd_data[21]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[21]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_10 
       (.I0(tagged_frame_transed_reg[21]),
        .I1(frame_1024_max_transed_reg[21]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[21]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[21]),
        .O(\stat_rd_data[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_11 
       (.I0(multicast_received_good_reg[21]),
        .I1(broadcast_received_good_reg[21]),
        .I2(out[1]),
        .I3(fcs_error_reg[21]),
        .I4(out[0]),
        .I5(frame_received_good_reg[21]),
        .O(\stat_rd_data[21]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_12 
       (.I0(frame_256_511_good_reg[21]),
        .I1(frame_128_255_good_reg[21]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[21]),
        .I4(out[0]),
        .I5(frame_64_good_reg[21]),
        .O(\stat_rd_data[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_13 
       (.I0(lt_out_range_reg[21]),
        .I1(control_frame_good_reg[21]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[21]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[21]),
        .O(\stat_rd_data[21]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_14 
       (.I0(oversize_frame_good_reg[21]),
        .I1(unsupported_control_frame_reg[21]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[21]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[21]),
        .O(\stat_rd_data[21]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_2 
       (.I0(\stat_rd_data_reg[21]_i_4_n_0 ),
        .I1(\stat_rd_data[21]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[21]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[21]_i_7_n_0 ),
        .O(\stat_rd_data[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_3 
       (.I0(total_bytes_transed_reg[21]),
        .I1(total_bytes_recved_reg[21]),
        .I2(out[1]),
        .I3(fragment_frame_reg[21]),
        .I4(out[0]),
        .I5(undersize_frame_reg[21]),
        .O(\stat_rd_data[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[21]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[21]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[21]),
        .I5(pause_frame_transed_reg[21]),
        .O(\stat_rd_data[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_6 
       (.I0(frame_128_255_transed_reg[21]),
        .I1(frame_65_127_transed_reg[21]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[21]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[21]),
        .O(\stat_rd_data[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[21]_i_7 
       (.I0(underrun_error_reg[21]),
        .I1(multicast_frame_transed_reg[21]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[21]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[21]),
        .O(\stat_rd_data[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[22]_i_1 
       (.I0(\stat_rd_data[22]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[22]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[22]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_10 
       (.I0(tagged_frame_transed_reg[22]),
        .I1(frame_1024_max_transed_reg[22]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[22]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[22]),
        .O(\stat_rd_data[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_11 
       (.I0(multicast_received_good_reg[22]),
        .I1(broadcast_received_good_reg[22]),
        .I2(out[1]),
        .I3(fcs_error_reg[22]),
        .I4(out[0]),
        .I5(frame_received_good_reg[22]),
        .O(\stat_rd_data[22]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_12 
       (.I0(frame_256_511_good_reg[22]),
        .I1(frame_128_255_good_reg[22]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[22]),
        .I4(out[0]),
        .I5(frame_64_good_reg[22]),
        .O(\stat_rd_data[22]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_13 
       (.I0(lt_out_range_reg[22]),
        .I1(control_frame_good_reg[22]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[22]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[22]),
        .O(\stat_rd_data[22]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_14 
       (.I0(oversize_frame_good_reg[22]),
        .I1(unsupported_control_frame_reg[22]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[22]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[22]),
        .O(\stat_rd_data[22]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_2 
       (.I0(\stat_rd_data_reg[22]_i_4_n_0 ),
        .I1(\stat_rd_data[22]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[22]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[22]_i_7_n_0 ),
        .O(\stat_rd_data[22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_3 
       (.I0(total_bytes_transed_reg[22]),
        .I1(total_bytes_recved_reg[22]),
        .I2(out[1]),
        .I3(fragment_frame_reg[22]),
        .I4(out[0]),
        .I5(undersize_frame_reg[22]),
        .O(\stat_rd_data[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[22]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[22]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[22]),
        .I5(pause_frame_transed_reg[22]),
        .O(\stat_rd_data[22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_6 
       (.I0(frame_128_255_transed_reg[22]),
        .I1(frame_65_127_transed_reg[22]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[22]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[22]),
        .O(\stat_rd_data[22]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[22]_i_7 
       (.I0(underrun_error_reg[22]),
        .I1(multicast_frame_transed_reg[22]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[22]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[22]),
        .O(\stat_rd_data[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[23]_i_1 
       (.I0(\stat_rd_data[23]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[23]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_10 
       (.I0(tagged_frame_transed_reg[23]),
        .I1(frame_1024_max_transed_reg[23]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[23]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[23]),
        .O(\stat_rd_data[23]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_11 
       (.I0(multicast_received_good_reg[23]),
        .I1(broadcast_received_good_reg[23]),
        .I2(out[1]),
        .I3(fcs_error_reg[23]),
        .I4(out[0]),
        .I5(frame_received_good_reg[23]),
        .O(\stat_rd_data[23]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_12 
       (.I0(frame_256_511_good_reg[23]),
        .I1(frame_128_255_good_reg[23]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[23]),
        .I4(out[0]),
        .I5(frame_64_good_reg[23]),
        .O(\stat_rd_data[23]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_13 
       (.I0(lt_out_range_reg[23]),
        .I1(control_frame_good_reg[23]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[23]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[23]),
        .O(\stat_rd_data[23]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_14 
       (.I0(oversize_frame_good_reg[23]),
        .I1(unsupported_control_frame_reg[23]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[23]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[23]),
        .O(\stat_rd_data[23]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_2 
       (.I0(\stat_rd_data_reg[23]_i_4_n_0 ),
        .I1(\stat_rd_data[23]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[23]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[23]_i_7_n_0 ),
        .O(\stat_rd_data[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_3 
       (.I0(total_bytes_transed_reg[23]),
        .I1(total_bytes_recved_reg[23]),
        .I2(out[1]),
        .I3(fragment_frame_reg[23]),
        .I4(out[0]),
        .I5(undersize_frame_reg[23]),
        .O(\stat_rd_data[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[23]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[23]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[23]),
        .I5(pause_frame_transed_reg[23]),
        .O(\stat_rd_data[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_6 
       (.I0(frame_128_255_transed_reg[23]),
        .I1(frame_65_127_transed_reg[23]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[23]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[23]),
        .O(\stat_rd_data[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[23]_i_7 
       (.I0(underrun_error_reg[23]),
        .I1(multicast_frame_transed_reg[23]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[23]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[23]),
        .O(\stat_rd_data[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[24]_i_1 
       (.I0(\stat_rd_data[24]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[24]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_10 
       (.I0(tagged_frame_transed_reg[24]),
        .I1(frame_1024_max_transed_reg[24]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[24]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[24]),
        .O(\stat_rd_data[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_11 
       (.I0(multicast_received_good_reg[24]),
        .I1(broadcast_received_good_reg[24]),
        .I2(out[1]),
        .I3(fcs_error_reg[24]),
        .I4(out[0]),
        .I5(frame_received_good_reg[24]),
        .O(\stat_rd_data[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_12 
       (.I0(frame_256_511_good_reg[24]),
        .I1(frame_128_255_good_reg[24]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[24]),
        .I4(out[0]),
        .I5(frame_64_good_reg[24]),
        .O(\stat_rd_data[24]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_13 
       (.I0(lt_out_range_reg[24]),
        .I1(control_frame_good_reg[24]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[24]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[24]),
        .O(\stat_rd_data[24]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_14 
       (.I0(oversize_frame_good_reg[24]),
        .I1(unsupported_control_frame_reg[24]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[24]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[24]),
        .O(\stat_rd_data[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_2 
       (.I0(\stat_rd_data_reg[24]_i_4_n_0 ),
        .I1(\stat_rd_data[24]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[24]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[24]_i_7_n_0 ),
        .O(\stat_rd_data[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_3 
       (.I0(total_bytes_transed_reg[24]),
        .I1(total_bytes_recved_reg[24]),
        .I2(out[1]),
        .I3(fragment_frame_reg[24]),
        .I4(out[0]),
        .I5(undersize_frame_reg[24]),
        .O(\stat_rd_data[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[24]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[24]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[24]),
        .I5(pause_frame_transed_reg[24]),
        .O(\stat_rd_data[24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_6 
       (.I0(frame_128_255_transed_reg[24]),
        .I1(frame_65_127_transed_reg[24]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[24]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[24]),
        .O(\stat_rd_data[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[24]_i_7 
       (.I0(underrun_error_reg[24]),
        .I1(multicast_frame_transed_reg[24]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[24]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[24]),
        .O(\stat_rd_data[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[25]_i_1 
       (.I0(\stat_rd_data[25]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[25]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_10 
       (.I0(tagged_frame_transed_reg[25]),
        .I1(frame_1024_max_transed_reg[25]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[25]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[25]),
        .O(\stat_rd_data[25]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_11 
       (.I0(multicast_received_good_reg[25]),
        .I1(broadcast_received_good_reg[25]),
        .I2(out[1]),
        .I3(fcs_error_reg[25]),
        .I4(out[0]),
        .I5(frame_received_good_reg[25]),
        .O(\stat_rd_data[25]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_12 
       (.I0(frame_256_511_good_reg[25]),
        .I1(frame_128_255_good_reg[25]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[25]),
        .I4(out[0]),
        .I5(frame_64_good_reg[25]),
        .O(\stat_rd_data[25]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_13 
       (.I0(lt_out_range_reg[25]),
        .I1(control_frame_good_reg[25]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[25]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[25]),
        .O(\stat_rd_data[25]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_14 
       (.I0(oversize_frame_good_reg[25]),
        .I1(unsupported_control_frame_reg[25]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[25]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[25]),
        .O(\stat_rd_data[25]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_2 
       (.I0(\stat_rd_data_reg[25]_i_4_n_0 ),
        .I1(\stat_rd_data[25]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[25]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[25]_i_7_n_0 ),
        .O(\stat_rd_data[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_3 
       (.I0(total_bytes_transed_reg[25]),
        .I1(total_bytes_recved_reg[25]),
        .I2(out[1]),
        .I3(fragment_frame_reg[25]),
        .I4(out[0]),
        .I5(undersize_frame_reg[25]),
        .O(\stat_rd_data[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[25]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[25]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[25]),
        .I5(pause_frame_transed_reg[25]),
        .O(\stat_rd_data[25]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_6 
       (.I0(frame_128_255_transed_reg[25]),
        .I1(frame_65_127_transed_reg[25]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[25]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[25]),
        .O(\stat_rd_data[25]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[25]_i_7 
       (.I0(underrun_error_reg[25]),
        .I1(multicast_frame_transed_reg[25]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[25]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[25]),
        .O(\stat_rd_data[25]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[26]_i_1 
       (.I0(\stat_rd_data[26]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[26]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[26]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_10 
       (.I0(tagged_frame_transed_reg[26]),
        .I1(frame_1024_max_transed_reg[26]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[26]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[26]),
        .O(\stat_rd_data[26]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_11 
       (.I0(multicast_received_good_reg[26]),
        .I1(broadcast_received_good_reg[26]),
        .I2(out[1]),
        .I3(fcs_error_reg[26]),
        .I4(out[0]),
        .I5(frame_received_good_reg[26]),
        .O(\stat_rd_data[26]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_12 
       (.I0(frame_256_511_good_reg[26]),
        .I1(frame_128_255_good_reg[26]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[26]),
        .I4(out[0]),
        .I5(frame_64_good_reg[26]),
        .O(\stat_rd_data[26]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_13 
       (.I0(lt_out_range_reg[26]),
        .I1(control_frame_good_reg[26]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[26]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[26]),
        .O(\stat_rd_data[26]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_14 
       (.I0(oversize_frame_good_reg[26]),
        .I1(unsupported_control_frame_reg[26]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[26]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[26]),
        .O(\stat_rd_data[26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_2 
       (.I0(\stat_rd_data_reg[26]_i_4_n_0 ),
        .I1(\stat_rd_data[26]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[26]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[26]_i_7_n_0 ),
        .O(\stat_rd_data[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_3 
       (.I0(total_bytes_transed_reg[26]),
        .I1(total_bytes_recved_reg[26]),
        .I2(out[1]),
        .I3(fragment_frame_reg[26]),
        .I4(out[0]),
        .I5(undersize_frame_reg[26]),
        .O(\stat_rd_data[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[26]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[26]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[26]),
        .I5(pause_frame_transed_reg[26]),
        .O(\stat_rd_data[26]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_6 
       (.I0(frame_128_255_transed_reg[26]),
        .I1(frame_65_127_transed_reg[26]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[26]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[26]),
        .O(\stat_rd_data[26]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[26]_i_7 
       (.I0(underrun_error_reg[26]),
        .I1(multicast_frame_transed_reg[26]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[26]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[26]),
        .O(\stat_rd_data[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[27]_i_1 
       (.I0(\stat_rd_data[27]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[27]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[27]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_10 
       (.I0(tagged_frame_transed_reg[27]),
        .I1(frame_1024_max_transed_reg[27]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[27]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[27]),
        .O(\stat_rd_data[27]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_11 
       (.I0(multicast_received_good_reg[27]),
        .I1(broadcast_received_good_reg[27]),
        .I2(out[1]),
        .I3(fcs_error_reg[27]),
        .I4(out[0]),
        .I5(frame_received_good_reg[27]),
        .O(\stat_rd_data[27]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_12 
       (.I0(frame_256_511_good_reg[27]),
        .I1(frame_128_255_good_reg[27]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[27]),
        .I4(out[0]),
        .I5(frame_64_good_reg[27]),
        .O(\stat_rd_data[27]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_13 
       (.I0(lt_out_range_reg[27]),
        .I1(control_frame_good_reg[27]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[27]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[27]),
        .O(\stat_rd_data[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_14 
       (.I0(oversize_frame_good_reg[27]),
        .I1(unsupported_control_frame_reg[27]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[27]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[27]),
        .O(\stat_rd_data[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_2 
       (.I0(\stat_rd_data_reg[27]_i_4_n_0 ),
        .I1(\stat_rd_data[27]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[27]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[27]_i_7_n_0 ),
        .O(\stat_rd_data[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_3 
       (.I0(total_bytes_transed_reg[27]),
        .I1(total_bytes_recved_reg[27]),
        .I2(out[1]),
        .I3(fragment_frame_reg[27]),
        .I4(out[0]),
        .I5(undersize_frame_reg[27]),
        .O(\stat_rd_data[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[27]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[27]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[27]),
        .I5(pause_frame_transed_reg[27]),
        .O(\stat_rd_data[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_6 
       (.I0(frame_128_255_transed_reg[27]),
        .I1(frame_65_127_transed_reg[27]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[27]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[27]),
        .O(\stat_rd_data[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[27]_i_7 
       (.I0(underrun_error_reg[27]),
        .I1(multicast_frame_transed_reg[27]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[27]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[27]),
        .O(\stat_rd_data[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[28]_i_1 
       (.I0(\stat_rd_data[28]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[28]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_10 
       (.I0(tagged_frame_transed_reg[28]),
        .I1(frame_1024_max_transed_reg[28]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[28]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[28]),
        .O(\stat_rd_data[28]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_11 
       (.I0(multicast_received_good_reg[28]),
        .I1(broadcast_received_good_reg[28]),
        .I2(out[1]),
        .I3(fcs_error_reg[28]),
        .I4(out[0]),
        .I5(frame_received_good_reg[28]),
        .O(\stat_rd_data[28]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_12 
       (.I0(frame_256_511_good_reg[28]),
        .I1(frame_128_255_good_reg[28]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[28]),
        .I4(out[0]),
        .I5(frame_64_good_reg[28]),
        .O(\stat_rd_data[28]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_13 
       (.I0(lt_out_range_reg[28]),
        .I1(control_frame_good_reg[28]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[28]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[28]),
        .O(\stat_rd_data[28]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_14 
       (.I0(oversize_frame_good_reg[28]),
        .I1(unsupported_control_frame_reg[28]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[28]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[28]),
        .O(\stat_rd_data[28]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_2 
       (.I0(\stat_rd_data_reg[28]_i_4_n_0 ),
        .I1(\stat_rd_data[28]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[28]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[28]_i_7_n_0 ),
        .O(\stat_rd_data[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_3 
       (.I0(total_bytes_transed_reg[28]),
        .I1(total_bytes_recved_reg[28]),
        .I2(out[1]),
        .I3(fragment_frame_reg[28]),
        .I4(out[0]),
        .I5(undersize_frame_reg[28]),
        .O(\stat_rd_data[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[28]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[28]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[28]),
        .I5(pause_frame_transed_reg[28]),
        .O(\stat_rd_data[28]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_6 
       (.I0(frame_128_255_transed_reg[28]),
        .I1(frame_65_127_transed_reg[28]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[28]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[28]),
        .O(\stat_rd_data[28]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[28]_i_7 
       (.I0(underrun_error_reg[28]),
        .I1(multicast_frame_transed_reg[28]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[28]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[28]),
        .O(\stat_rd_data[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[29]_i_1 
       (.I0(\stat_rd_data[29]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[29]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_10 
       (.I0(tagged_frame_transed_reg[29]),
        .I1(frame_1024_max_transed_reg[29]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[29]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[29]),
        .O(\stat_rd_data[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_11 
       (.I0(multicast_received_good_reg[29]),
        .I1(broadcast_received_good_reg[29]),
        .I2(out[1]),
        .I3(fcs_error_reg[29]),
        .I4(out[0]),
        .I5(frame_received_good_reg[29]),
        .O(\stat_rd_data[29]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_12 
       (.I0(frame_256_511_good_reg[29]),
        .I1(frame_128_255_good_reg[29]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[29]),
        .I4(out[0]),
        .I5(frame_64_good_reg[29]),
        .O(\stat_rd_data[29]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_13 
       (.I0(lt_out_range_reg[29]),
        .I1(control_frame_good_reg[29]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[29]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[29]),
        .O(\stat_rd_data[29]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_14 
       (.I0(oversize_frame_good_reg[29]),
        .I1(unsupported_control_frame_reg[29]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[29]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[29]),
        .O(\stat_rd_data[29]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_2 
       (.I0(\stat_rd_data_reg[29]_i_4_n_0 ),
        .I1(\stat_rd_data[29]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[29]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[29]_i_7_n_0 ),
        .O(\stat_rd_data[29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_3 
       (.I0(total_bytes_transed_reg[29]),
        .I1(total_bytes_recved_reg[29]),
        .I2(out[1]),
        .I3(fragment_frame_reg[29]),
        .I4(out[0]),
        .I5(undersize_frame_reg[29]),
        .O(\stat_rd_data[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[29]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[29]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[29]),
        .I5(pause_frame_transed_reg[29]),
        .O(\stat_rd_data[29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_6 
       (.I0(frame_128_255_transed_reg[29]),
        .I1(frame_65_127_transed_reg[29]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[29]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[29]),
        .O(\stat_rd_data[29]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[29]_i_7 
       (.I0(underrun_error_reg[29]),
        .I1(multicast_frame_transed_reg[29]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[29]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[29]),
        .O(\stat_rd_data[29]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[2]_i_1 
       (.I0(\stat_rd_data[2]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[2]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_10 
       (.I0(tagged_frame_transed_reg[2]),
        .I1(frame_1024_max_transed_reg[2]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[2]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[2]),
        .O(\stat_rd_data[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_11 
       (.I0(multicast_received_good_reg[2]),
        .I1(broadcast_received_good_reg[2]),
        .I2(out[1]),
        .I3(fcs_error_reg[2]),
        .I4(out[0]),
        .I5(frame_received_good_reg[2]),
        .O(\stat_rd_data[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_12 
       (.I0(frame_256_511_good_reg[2]),
        .I1(frame_128_255_good_reg[2]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[2]),
        .I4(out[0]),
        .I5(frame_64_good_reg[2]),
        .O(\stat_rd_data[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_13 
       (.I0(lt_out_range_reg[2]),
        .I1(control_frame_good_reg[2]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[2]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[2]),
        .O(\stat_rd_data[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_14 
       (.I0(oversize_frame_good_reg[2]),
        .I1(unsupported_control_frame_reg[2]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[2]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[2]),
        .O(\stat_rd_data[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_2 
       (.I0(\stat_rd_data_reg[2]_i_4_n_0 ),
        .I1(\stat_rd_data[2]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[2]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[2]_i_7_n_0 ),
        .O(\stat_rd_data[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_3 
       (.I0(total_bytes_transed_reg[2]),
        .I1(total_bytes_recved_reg[2]),
        .I2(out[1]),
        .I3(fragment_frame_reg[2]),
        .I4(out[0]),
        .I5(undersize_frame_reg[2]),
        .O(\stat_rd_data[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[2]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[2]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[2]),
        .I5(pause_frame_transed_reg[2]),
        .O(\stat_rd_data[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_6 
       (.I0(frame_128_255_transed_reg[2]),
        .I1(frame_65_127_transed_reg[2]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[2]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[2]),
        .O(\stat_rd_data[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[2]_i_7 
       (.I0(underrun_error_reg[2]),
        .I1(multicast_frame_transed_reg[2]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[2]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[2]),
        .O(\stat_rd_data[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[30]_i_1 
       (.I0(\stat_rd_data[30]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[30]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_10 
       (.I0(tagged_frame_transed_reg[30]),
        .I1(frame_1024_max_transed_reg[30]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[30]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[30]),
        .O(\stat_rd_data[30]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_11 
       (.I0(multicast_received_good_reg[30]),
        .I1(broadcast_received_good_reg[30]),
        .I2(out[1]),
        .I3(fcs_error_reg[30]),
        .I4(out[0]),
        .I5(frame_received_good_reg[30]),
        .O(\stat_rd_data[30]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_12 
       (.I0(frame_256_511_good_reg[30]),
        .I1(frame_128_255_good_reg[30]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[30]),
        .I4(out[0]),
        .I5(frame_64_good_reg[30]),
        .O(\stat_rd_data[30]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_13 
       (.I0(lt_out_range_reg[30]),
        .I1(control_frame_good_reg[30]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[30]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[30]),
        .O(\stat_rd_data[30]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_14 
       (.I0(oversize_frame_good_reg[30]),
        .I1(unsupported_control_frame_reg[30]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[30]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[30]),
        .O(\stat_rd_data[30]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_2 
       (.I0(\stat_rd_data_reg[30]_i_4_n_0 ),
        .I1(\stat_rd_data[30]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[30]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[30]_i_7_n_0 ),
        .O(\stat_rd_data[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_3 
       (.I0(total_bytes_transed_reg[30]),
        .I1(total_bytes_recved_reg[30]),
        .I2(out[1]),
        .I3(fragment_frame_reg[30]),
        .I4(out[0]),
        .I5(undersize_frame_reg[30]),
        .O(\stat_rd_data[30]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[30]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[30]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[30]),
        .I5(pause_frame_transed_reg[30]),
        .O(\stat_rd_data[30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_6 
       (.I0(frame_128_255_transed_reg[30]),
        .I1(frame_65_127_transed_reg[30]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[30]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[30]),
        .O(\stat_rd_data[30]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[30]_i_7 
       (.I0(underrun_error_reg[30]),
        .I1(multicast_frame_transed_reg[30]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[30]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[30]),
        .O(\stat_rd_data[30]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[31]_i_1 
       (.I0(\stat_rd_data[31]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[31]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[31]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_10 
       (.I0(tagged_frame_transed_reg[31]),
        .I1(frame_1024_max_transed_reg[31]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[31]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[31]),
        .O(\stat_rd_data[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_11 
       (.I0(multicast_received_good_reg[31]),
        .I1(broadcast_received_good_reg[31]),
        .I2(out[1]),
        .I3(fcs_error_reg[31]),
        .I4(out[0]),
        .I5(frame_received_good_reg[31]),
        .O(\stat_rd_data[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_12 
       (.I0(frame_256_511_good_reg[31]),
        .I1(frame_128_255_good_reg[31]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[31]),
        .I4(out[0]),
        .I5(frame_64_good_reg[31]),
        .O(\stat_rd_data[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_13 
       (.I0(lt_out_range_reg[31]),
        .I1(control_frame_good_reg[31]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[31]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[31]),
        .O(\stat_rd_data[31]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_14 
       (.I0(oversize_frame_good_reg[31]),
        .I1(unsupported_control_frame_reg[31]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[31]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[31]),
        .O(\stat_rd_data[31]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_2 
       (.I0(\stat_rd_data_reg[31]_i_4_n_0 ),
        .I1(\stat_rd_data[31]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[31]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[31]_i_7_n_0 ),
        .O(\stat_rd_data[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_3 
       (.I0(total_bytes_transed_reg[31]),
        .I1(total_bytes_recved_reg[31]),
        .I2(out[1]),
        .I3(fragment_frame_reg[31]),
        .I4(out[0]),
        .I5(undersize_frame_reg[31]),
        .O(\stat_rd_data[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[31]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[31]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[31]),
        .I5(pause_frame_transed_reg[31]),
        .O(\stat_rd_data[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_6 
       (.I0(frame_128_255_transed_reg[31]),
        .I1(frame_65_127_transed_reg[31]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[31]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[31]),
        .O(\stat_rd_data[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[31]_i_7 
       (.I0(underrun_error_reg[31]),
        .I1(multicast_frame_transed_reg[31]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[31]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[31]),
        .O(\stat_rd_data[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[32]_i_1 
       (.I0(\stat_rd_data[32]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[32]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[32]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_10 
       (.I0(tagged_frame_transed_reg[32]),
        .I1(frame_1024_max_transed_reg[32]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[32]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[32]),
        .O(\stat_rd_data[32]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_11 
       (.I0(multicast_received_good_reg[32]),
        .I1(broadcast_received_good_reg[32]),
        .I2(out[1]),
        .I3(fcs_error_reg[32]),
        .I4(out[0]),
        .I5(frame_received_good_reg[32]),
        .O(\stat_rd_data[32]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_12 
       (.I0(frame_256_511_good_reg[32]),
        .I1(frame_128_255_good_reg[32]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[32]),
        .I4(out[0]),
        .I5(frame_64_good_reg[32]),
        .O(\stat_rd_data[32]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_13 
       (.I0(lt_out_range_reg[32]),
        .I1(control_frame_good_reg[32]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[32]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[32]),
        .O(\stat_rd_data[32]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_14 
       (.I0(oversize_frame_good_reg[32]),
        .I1(unsupported_control_frame_reg[32]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[32]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[32]),
        .O(\stat_rd_data[32]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_2 
       (.I0(\stat_rd_data_reg[32]_i_4_n_0 ),
        .I1(\stat_rd_data[32]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[32]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[32]_i_7_n_0 ),
        .O(\stat_rd_data[32]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_3 
       (.I0(total_bytes_transed_reg[32]),
        .I1(total_bytes_recved_reg[32]),
        .I2(out[1]),
        .I3(fragment_frame_reg[32]),
        .I4(out[0]),
        .I5(undersize_frame_reg[32]),
        .O(\stat_rd_data[32]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[32]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[32]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[32]),
        .I5(pause_frame_transed_reg[32]),
        .O(\stat_rd_data[32]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_6 
       (.I0(frame_128_255_transed_reg[32]),
        .I1(frame_65_127_transed_reg[32]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[32]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[32]),
        .O(\stat_rd_data[32]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[32]_i_7 
       (.I0(underrun_error_reg[32]),
        .I1(multicast_frame_transed_reg[32]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[32]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[32]),
        .O(\stat_rd_data[32]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[33]_i_1 
       (.I0(\stat_rd_data[33]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[33]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[33]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_10 
       (.I0(tagged_frame_transed_reg[33]),
        .I1(frame_1024_max_transed_reg[33]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[33]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[33]),
        .O(\stat_rd_data[33]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_11 
       (.I0(multicast_received_good_reg[33]),
        .I1(broadcast_received_good_reg[33]),
        .I2(out[1]),
        .I3(fcs_error_reg[33]),
        .I4(out[0]),
        .I5(frame_received_good_reg[33]),
        .O(\stat_rd_data[33]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_12 
       (.I0(frame_256_511_good_reg[33]),
        .I1(frame_128_255_good_reg[33]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[33]),
        .I4(out[0]),
        .I5(frame_64_good_reg[33]),
        .O(\stat_rd_data[33]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_13 
       (.I0(lt_out_range_reg[33]),
        .I1(control_frame_good_reg[33]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[33]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[33]),
        .O(\stat_rd_data[33]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_14 
       (.I0(oversize_frame_good_reg[33]),
        .I1(unsupported_control_frame_reg[33]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[33]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[33]),
        .O(\stat_rd_data[33]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_2 
       (.I0(\stat_rd_data_reg[33]_i_4_n_0 ),
        .I1(\stat_rd_data[33]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[33]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[33]_i_7_n_0 ),
        .O(\stat_rd_data[33]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_3 
       (.I0(total_bytes_transed_reg[33]),
        .I1(total_bytes_recved_reg[33]),
        .I2(out[1]),
        .I3(fragment_frame_reg[33]),
        .I4(out[0]),
        .I5(undersize_frame_reg[33]),
        .O(\stat_rd_data[33]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[33]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[33]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[33]),
        .I5(pause_frame_transed_reg[33]),
        .O(\stat_rd_data[33]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_6 
       (.I0(frame_128_255_transed_reg[33]),
        .I1(frame_65_127_transed_reg[33]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[33]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[33]),
        .O(\stat_rd_data[33]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[33]_i_7 
       (.I0(underrun_error_reg[33]),
        .I1(multicast_frame_transed_reg[33]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[33]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[33]),
        .O(\stat_rd_data[33]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[34]_i_1 
       (.I0(\stat_rd_data[34]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[34]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[34]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_10 
       (.I0(tagged_frame_transed_reg[34]),
        .I1(frame_1024_max_transed_reg[34]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[34]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[34]),
        .O(\stat_rd_data[34]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_11 
       (.I0(multicast_received_good_reg[34]),
        .I1(broadcast_received_good_reg[34]),
        .I2(out[1]),
        .I3(fcs_error_reg[34]),
        .I4(out[0]),
        .I5(frame_received_good_reg[34]),
        .O(\stat_rd_data[34]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_12 
       (.I0(frame_256_511_good_reg[34]),
        .I1(frame_128_255_good_reg[34]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[34]),
        .I4(out[0]),
        .I5(frame_64_good_reg[34]),
        .O(\stat_rd_data[34]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_13 
       (.I0(lt_out_range_reg[34]),
        .I1(control_frame_good_reg[34]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[34]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[34]),
        .O(\stat_rd_data[34]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_14 
       (.I0(oversize_frame_good_reg[34]),
        .I1(unsupported_control_frame_reg[34]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[34]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[34]),
        .O(\stat_rd_data[34]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_2 
       (.I0(\stat_rd_data_reg[34]_i_4_n_0 ),
        .I1(\stat_rd_data[34]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[34]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[34]_i_7_n_0 ),
        .O(\stat_rd_data[34]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_3 
       (.I0(total_bytes_transed_reg[34]),
        .I1(total_bytes_recved_reg[34]),
        .I2(out[1]),
        .I3(fragment_frame_reg[34]),
        .I4(out[0]),
        .I5(undersize_frame_reg[34]),
        .O(\stat_rd_data[34]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[34]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[34]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[34]),
        .I5(pause_frame_transed_reg[34]),
        .O(\stat_rd_data[34]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_6 
       (.I0(frame_128_255_transed_reg[34]),
        .I1(frame_65_127_transed_reg[34]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[34]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[34]),
        .O(\stat_rd_data[34]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[34]_i_7 
       (.I0(underrun_error_reg[34]),
        .I1(multicast_frame_transed_reg[34]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[34]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[34]),
        .O(\stat_rd_data[34]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[35]_i_1 
       (.I0(\stat_rd_data[35]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[35]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[35]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_10 
       (.I0(tagged_frame_transed_reg[35]),
        .I1(frame_1024_max_transed_reg[35]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[35]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[35]),
        .O(\stat_rd_data[35]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_11 
       (.I0(multicast_received_good_reg[35]),
        .I1(broadcast_received_good_reg[35]),
        .I2(out[1]),
        .I3(fcs_error_reg[35]),
        .I4(out[0]),
        .I5(frame_received_good_reg[35]),
        .O(\stat_rd_data[35]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_12 
       (.I0(frame_256_511_good_reg[35]),
        .I1(frame_128_255_good_reg[35]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[35]),
        .I4(out[0]),
        .I5(frame_64_good_reg[35]),
        .O(\stat_rd_data[35]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_13 
       (.I0(lt_out_range_reg[35]),
        .I1(control_frame_good_reg[35]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[35]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[35]),
        .O(\stat_rd_data[35]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_14 
       (.I0(oversize_frame_good_reg[35]),
        .I1(unsupported_control_frame_reg[35]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[35]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[35]),
        .O(\stat_rd_data[35]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_2 
       (.I0(\stat_rd_data_reg[35]_i_4_n_0 ),
        .I1(\stat_rd_data[35]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[35]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[35]_i_7_n_0 ),
        .O(\stat_rd_data[35]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_3 
       (.I0(total_bytes_transed_reg[35]),
        .I1(total_bytes_recved_reg[35]),
        .I2(out[1]),
        .I3(fragment_frame_reg[35]),
        .I4(out[0]),
        .I5(undersize_frame_reg[35]),
        .O(\stat_rd_data[35]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[35]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[35]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[35]),
        .I5(pause_frame_transed_reg[35]),
        .O(\stat_rd_data[35]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_6 
       (.I0(frame_128_255_transed_reg[35]),
        .I1(frame_65_127_transed_reg[35]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[35]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[35]),
        .O(\stat_rd_data[35]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[35]_i_7 
       (.I0(underrun_error_reg[35]),
        .I1(multicast_frame_transed_reg[35]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[35]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[35]),
        .O(\stat_rd_data[35]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[36]_i_1 
       (.I0(\stat_rd_data[36]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[36]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[36]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_10 
       (.I0(tagged_frame_transed_reg[36]),
        .I1(frame_1024_max_transed_reg[36]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[36]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[36]),
        .O(\stat_rd_data[36]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_11 
       (.I0(multicast_received_good_reg[36]),
        .I1(broadcast_received_good_reg[36]),
        .I2(out[1]),
        .I3(fcs_error_reg[36]),
        .I4(out[0]),
        .I5(frame_received_good_reg[36]),
        .O(\stat_rd_data[36]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_12 
       (.I0(frame_256_511_good_reg[36]),
        .I1(frame_128_255_good_reg[36]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[36]),
        .I4(out[0]),
        .I5(frame_64_good_reg[36]),
        .O(\stat_rd_data[36]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_13 
       (.I0(lt_out_range_reg[36]),
        .I1(control_frame_good_reg[36]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[36]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[36]),
        .O(\stat_rd_data[36]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_14 
       (.I0(oversize_frame_good_reg[36]),
        .I1(unsupported_control_frame_reg[36]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[36]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[36]),
        .O(\stat_rd_data[36]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_2 
       (.I0(\stat_rd_data_reg[36]_i_4_n_0 ),
        .I1(\stat_rd_data[36]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[36]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[36]_i_7_n_0 ),
        .O(\stat_rd_data[36]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_3 
       (.I0(total_bytes_transed_reg[36]),
        .I1(total_bytes_recved_reg[36]),
        .I2(out[1]),
        .I3(fragment_frame_reg[36]),
        .I4(out[0]),
        .I5(undersize_frame_reg[36]),
        .O(\stat_rd_data[36]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[36]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[36]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[36]),
        .I5(pause_frame_transed_reg[36]),
        .O(\stat_rd_data[36]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_6 
       (.I0(frame_128_255_transed_reg[36]),
        .I1(frame_65_127_transed_reg[36]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[36]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[36]),
        .O(\stat_rd_data[36]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[36]_i_7 
       (.I0(underrun_error_reg[36]),
        .I1(multicast_frame_transed_reg[36]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[36]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[36]),
        .O(\stat_rd_data[36]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[37]_i_1 
       (.I0(\stat_rd_data[37]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[37]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[37]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_10 
       (.I0(tagged_frame_transed_reg[37]),
        .I1(frame_1024_max_transed_reg[37]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[37]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[37]),
        .O(\stat_rd_data[37]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_11 
       (.I0(multicast_received_good_reg[37]),
        .I1(broadcast_received_good_reg[37]),
        .I2(out[1]),
        .I3(fcs_error_reg[37]),
        .I4(out[0]),
        .I5(frame_received_good_reg[37]),
        .O(\stat_rd_data[37]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_12 
       (.I0(frame_256_511_good_reg[37]),
        .I1(frame_128_255_good_reg[37]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[37]),
        .I4(out[0]),
        .I5(frame_64_good_reg[37]),
        .O(\stat_rd_data[37]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_13 
       (.I0(lt_out_range_reg[37]),
        .I1(control_frame_good_reg[37]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[37]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[37]),
        .O(\stat_rd_data[37]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_14 
       (.I0(oversize_frame_good_reg[37]),
        .I1(unsupported_control_frame_reg[37]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[37]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[37]),
        .O(\stat_rd_data[37]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_2 
       (.I0(\stat_rd_data_reg[37]_i_4_n_0 ),
        .I1(\stat_rd_data[37]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[37]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[37]_i_7_n_0 ),
        .O(\stat_rd_data[37]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_3 
       (.I0(total_bytes_transed_reg[37]),
        .I1(total_bytes_recved_reg[37]),
        .I2(out[1]),
        .I3(fragment_frame_reg[37]),
        .I4(out[0]),
        .I5(undersize_frame_reg[37]),
        .O(\stat_rd_data[37]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[37]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[37]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[37]),
        .I5(pause_frame_transed_reg[37]),
        .O(\stat_rd_data[37]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_6 
       (.I0(frame_128_255_transed_reg[37]),
        .I1(frame_65_127_transed_reg[37]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[37]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[37]),
        .O(\stat_rd_data[37]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[37]_i_7 
       (.I0(underrun_error_reg[37]),
        .I1(multicast_frame_transed_reg[37]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[37]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[37]),
        .O(\stat_rd_data[37]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[38]_i_1 
       (.I0(\stat_rd_data[38]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[38]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[38]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_10 
       (.I0(tagged_frame_transed_reg[38]),
        .I1(frame_1024_max_transed_reg[38]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[38]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[38]),
        .O(\stat_rd_data[38]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_11 
       (.I0(multicast_received_good_reg[38]),
        .I1(broadcast_received_good_reg[38]),
        .I2(out[1]),
        .I3(fcs_error_reg[38]),
        .I4(out[0]),
        .I5(frame_received_good_reg[38]),
        .O(\stat_rd_data[38]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_12 
       (.I0(frame_256_511_good_reg[38]),
        .I1(frame_128_255_good_reg[38]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[38]),
        .I4(out[0]),
        .I5(frame_64_good_reg[38]),
        .O(\stat_rd_data[38]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_13 
       (.I0(lt_out_range_reg[38]),
        .I1(control_frame_good_reg[38]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[38]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[38]),
        .O(\stat_rd_data[38]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_14 
       (.I0(oversize_frame_good_reg[38]),
        .I1(unsupported_control_frame_reg[38]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[38]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[38]),
        .O(\stat_rd_data[38]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_2 
       (.I0(\stat_rd_data_reg[38]_i_4_n_0 ),
        .I1(\stat_rd_data[38]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[38]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[38]_i_7_n_0 ),
        .O(\stat_rd_data[38]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_3 
       (.I0(total_bytes_transed_reg[38]),
        .I1(total_bytes_recved_reg[38]),
        .I2(out[1]),
        .I3(fragment_frame_reg[38]),
        .I4(out[0]),
        .I5(undersize_frame_reg[38]),
        .O(\stat_rd_data[38]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[38]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[38]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[38]),
        .I5(pause_frame_transed_reg[38]),
        .O(\stat_rd_data[38]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_6 
       (.I0(frame_128_255_transed_reg[38]),
        .I1(frame_65_127_transed_reg[38]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[38]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[38]),
        .O(\stat_rd_data[38]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[38]_i_7 
       (.I0(underrun_error_reg[38]),
        .I1(multicast_frame_transed_reg[38]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[38]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[38]),
        .O(\stat_rd_data[38]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[39]_i_1 
       (.I0(\stat_rd_data[39]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[39]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[39]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_10 
       (.I0(tagged_frame_transed_reg[39]),
        .I1(frame_1024_max_transed_reg[39]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[39]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[39]),
        .O(\stat_rd_data[39]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_11 
       (.I0(multicast_received_good_reg[39]),
        .I1(broadcast_received_good_reg[39]),
        .I2(out[1]),
        .I3(fcs_error_reg[39]),
        .I4(out[0]),
        .I5(frame_received_good_reg[39]),
        .O(\stat_rd_data[39]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_12 
       (.I0(frame_256_511_good_reg[39]),
        .I1(frame_128_255_good_reg[39]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[39]),
        .I4(out[0]),
        .I5(frame_64_good_reg[39]),
        .O(\stat_rd_data[39]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_13 
       (.I0(lt_out_range_reg[39]),
        .I1(control_frame_good_reg[39]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[39]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[39]),
        .O(\stat_rd_data[39]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_14 
       (.I0(oversize_frame_good_reg[39]),
        .I1(unsupported_control_frame_reg[39]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[39]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[39]),
        .O(\stat_rd_data[39]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_2 
       (.I0(\stat_rd_data_reg[39]_i_4_n_0 ),
        .I1(\stat_rd_data[39]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[39]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[39]_i_7_n_0 ),
        .O(\stat_rd_data[39]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_3 
       (.I0(total_bytes_transed_reg[39]),
        .I1(total_bytes_recved_reg[39]),
        .I2(out[1]),
        .I3(fragment_frame_reg[39]),
        .I4(out[0]),
        .I5(undersize_frame_reg[39]),
        .O(\stat_rd_data[39]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[39]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[39]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[39]),
        .I5(pause_frame_transed_reg[39]),
        .O(\stat_rd_data[39]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_6 
       (.I0(frame_128_255_transed_reg[39]),
        .I1(frame_65_127_transed_reg[39]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[39]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[39]),
        .O(\stat_rd_data[39]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[39]_i_7 
       (.I0(underrun_error_reg[39]),
        .I1(multicast_frame_transed_reg[39]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[39]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[39]),
        .O(\stat_rd_data[39]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[3]_i_1 
       (.I0(\stat_rd_data[3]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[3]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_10 
       (.I0(tagged_frame_transed_reg[3]),
        .I1(frame_1024_max_transed_reg[3]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[3]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[3]),
        .O(\stat_rd_data[3]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_11 
       (.I0(multicast_received_good_reg[3]),
        .I1(broadcast_received_good_reg[3]),
        .I2(out[1]),
        .I3(fcs_error_reg[3]),
        .I4(out[0]),
        .I5(frame_received_good_reg[3]),
        .O(\stat_rd_data[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_12 
       (.I0(frame_256_511_good_reg[3]),
        .I1(frame_128_255_good_reg[3]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[3]),
        .I4(out[0]),
        .I5(frame_64_good_reg[3]),
        .O(\stat_rd_data[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_13 
       (.I0(lt_out_range_reg[3]),
        .I1(control_frame_good_reg[3]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[3]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[3]),
        .O(\stat_rd_data[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_14 
       (.I0(oversize_frame_good_reg[3]),
        .I1(unsupported_control_frame_reg[3]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[3]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[3]),
        .O(\stat_rd_data[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_2 
       (.I0(\stat_rd_data_reg[3]_i_4_n_0 ),
        .I1(\stat_rd_data[3]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[3]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[3]_i_7_n_0 ),
        .O(\stat_rd_data[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_3 
       (.I0(total_bytes_transed_reg[3]),
        .I1(total_bytes_recved_reg[3]),
        .I2(out[1]),
        .I3(fragment_frame_reg[3]),
        .I4(out[0]),
        .I5(undersize_frame_reg[3]),
        .O(\stat_rd_data[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[3]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[3]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[3]),
        .I5(pause_frame_transed_reg[3]),
        .O(\stat_rd_data[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_6 
       (.I0(frame_128_255_transed_reg[3]),
        .I1(frame_65_127_transed_reg[3]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[3]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[3]),
        .O(\stat_rd_data[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[3]_i_7 
       (.I0(underrun_error_reg[3]),
        .I1(multicast_frame_transed_reg[3]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[3]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[3]),
        .O(\stat_rd_data[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[40]_i_1 
       (.I0(\stat_rd_data[40]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[40]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[40]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_10 
       (.I0(tagged_frame_transed_reg[40]),
        .I1(frame_1024_max_transed_reg[40]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[40]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[40]),
        .O(\stat_rd_data[40]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_11 
       (.I0(multicast_received_good_reg[40]),
        .I1(broadcast_received_good_reg[40]),
        .I2(out[1]),
        .I3(fcs_error_reg[40]),
        .I4(out[0]),
        .I5(frame_received_good_reg[40]),
        .O(\stat_rd_data[40]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_12 
       (.I0(frame_256_511_good_reg[40]),
        .I1(frame_128_255_good_reg[40]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[40]),
        .I4(out[0]),
        .I5(frame_64_good_reg[40]),
        .O(\stat_rd_data[40]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_13 
       (.I0(lt_out_range_reg[40]),
        .I1(control_frame_good_reg[40]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[40]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[40]),
        .O(\stat_rd_data[40]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_14 
       (.I0(oversize_frame_good_reg[40]),
        .I1(unsupported_control_frame_reg[40]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[40]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[40]),
        .O(\stat_rd_data[40]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_2 
       (.I0(\stat_rd_data_reg[40]_i_4_n_0 ),
        .I1(\stat_rd_data[40]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[40]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[40]_i_7_n_0 ),
        .O(\stat_rd_data[40]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_3 
       (.I0(total_bytes_transed_reg[40]),
        .I1(total_bytes_recved_reg[40]),
        .I2(out[1]),
        .I3(fragment_frame_reg[40]),
        .I4(out[0]),
        .I5(undersize_frame_reg[40]),
        .O(\stat_rd_data[40]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[40]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[40]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[40]),
        .I5(pause_frame_transed_reg[40]),
        .O(\stat_rd_data[40]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_6 
       (.I0(frame_128_255_transed_reg[40]),
        .I1(frame_65_127_transed_reg[40]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[40]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[40]),
        .O(\stat_rd_data[40]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[40]_i_7 
       (.I0(underrun_error_reg[40]),
        .I1(multicast_frame_transed_reg[40]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[40]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[40]),
        .O(\stat_rd_data[40]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[41]_i_1 
       (.I0(\stat_rd_data[41]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[41]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[41]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_10 
       (.I0(tagged_frame_transed_reg[41]),
        .I1(frame_1024_max_transed_reg[41]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[41]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[41]),
        .O(\stat_rd_data[41]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_11 
       (.I0(multicast_received_good_reg[41]),
        .I1(broadcast_received_good_reg[41]),
        .I2(out[1]),
        .I3(fcs_error_reg[41]),
        .I4(out[0]),
        .I5(frame_received_good_reg[41]),
        .O(\stat_rd_data[41]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_12 
       (.I0(frame_256_511_good_reg[41]),
        .I1(frame_128_255_good_reg[41]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[41]),
        .I4(out[0]),
        .I5(frame_64_good_reg[41]),
        .O(\stat_rd_data[41]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_13 
       (.I0(lt_out_range_reg[41]),
        .I1(control_frame_good_reg[41]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[41]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[41]),
        .O(\stat_rd_data[41]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_14 
       (.I0(oversize_frame_good_reg[41]),
        .I1(unsupported_control_frame_reg[41]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[41]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[41]),
        .O(\stat_rd_data[41]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_2 
       (.I0(\stat_rd_data_reg[41]_i_4_n_0 ),
        .I1(\stat_rd_data[41]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[41]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[41]_i_7_n_0 ),
        .O(\stat_rd_data[41]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_3 
       (.I0(total_bytes_transed_reg[41]),
        .I1(total_bytes_recved_reg[41]),
        .I2(out[1]),
        .I3(fragment_frame_reg[41]),
        .I4(out[0]),
        .I5(undersize_frame_reg[41]),
        .O(\stat_rd_data[41]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[41]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[41]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[41]),
        .I5(pause_frame_transed_reg[41]),
        .O(\stat_rd_data[41]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_6 
       (.I0(frame_128_255_transed_reg[41]),
        .I1(frame_65_127_transed_reg[41]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[41]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[41]),
        .O(\stat_rd_data[41]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[41]_i_7 
       (.I0(underrun_error_reg[41]),
        .I1(multicast_frame_transed_reg[41]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[41]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[41]),
        .O(\stat_rd_data[41]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[42]_i_1 
       (.I0(\stat_rd_data[42]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[42]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[42]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_10 
       (.I0(tagged_frame_transed_reg[42]),
        .I1(frame_1024_max_transed_reg[42]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[42]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[42]),
        .O(\stat_rd_data[42]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_11 
       (.I0(multicast_received_good_reg[42]),
        .I1(broadcast_received_good_reg[42]),
        .I2(out[1]),
        .I3(fcs_error_reg[42]),
        .I4(out[0]),
        .I5(frame_received_good_reg[42]),
        .O(\stat_rd_data[42]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_12 
       (.I0(frame_256_511_good_reg[42]),
        .I1(frame_128_255_good_reg[42]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[42]),
        .I4(out[0]),
        .I5(frame_64_good_reg[42]),
        .O(\stat_rd_data[42]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_13 
       (.I0(lt_out_range_reg[42]),
        .I1(control_frame_good_reg[42]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[42]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[42]),
        .O(\stat_rd_data[42]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_14 
       (.I0(oversize_frame_good_reg[42]),
        .I1(unsupported_control_frame_reg[42]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[42]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[42]),
        .O(\stat_rd_data[42]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_2 
       (.I0(\stat_rd_data_reg[42]_i_4_n_0 ),
        .I1(\stat_rd_data[42]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[42]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[42]_i_7_n_0 ),
        .O(\stat_rd_data[42]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_3 
       (.I0(total_bytes_transed_reg[42]),
        .I1(total_bytes_recved_reg[42]),
        .I2(out[1]),
        .I3(fragment_frame_reg[42]),
        .I4(out[0]),
        .I5(undersize_frame_reg[42]),
        .O(\stat_rd_data[42]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[42]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[42]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[42]),
        .I5(pause_frame_transed_reg[42]),
        .O(\stat_rd_data[42]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_6 
       (.I0(frame_128_255_transed_reg[42]),
        .I1(frame_65_127_transed_reg[42]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[42]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[42]),
        .O(\stat_rd_data[42]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[42]_i_7 
       (.I0(underrun_error_reg[42]),
        .I1(multicast_frame_transed_reg[42]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[42]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[42]),
        .O(\stat_rd_data[42]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[43]_i_1 
       (.I0(\stat_rd_data[43]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[43]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[43]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_10 
       (.I0(tagged_frame_transed_reg[43]),
        .I1(frame_1024_max_transed_reg[43]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[43]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[43]),
        .O(\stat_rd_data[43]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_11 
       (.I0(multicast_received_good_reg[43]),
        .I1(broadcast_received_good_reg[43]),
        .I2(out[1]),
        .I3(fcs_error_reg[43]),
        .I4(out[0]),
        .I5(frame_received_good_reg[43]),
        .O(\stat_rd_data[43]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_12 
       (.I0(frame_256_511_good_reg[43]),
        .I1(frame_128_255_good_reg[43]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[43]),
        .I4(out[0]),
        .I5(frame_64_good_reg[43]),
        .O(\stat_rd_data[43]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_13 
       (.I0(lt_out_range_reg[43]),
        .I1(control_frame_good_reg[43]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[43]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[43]),
        .O(\stat_rd_data[43]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_14 
       (.I0(oversize_frame_good_reg[43]),
        .I1(unsupported_control_frame_reg[43]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[43]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[43]),
        .O(\stat_rd_data[43]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_2 
       (.I0(\stat_rd_data_reg[43]_i_4_n_0 ),
        .I1(\stat_rd_data[43]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[43]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[43]_i_7_n_0 ),
        .O(\stat_rd_data[43]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_3 
       (.I0(total_bytes_transed_reg[43]),
        .I1(total_bytes_recved_reg[43]),
        .I2(out[1]),
        .I3(fragment_frame_reg[43]),
        .I4(out[0]),
        .I5(undersize_frame_reg[43]),
        .O(\stat_rd_data[43]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[43]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[43]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[43]),
        .I5(pause_frame_transed_reg[43]),
        .O(\stat_rd_data[43]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_6 
       (.I0(frame_128_255_transed_reg[43]),
        .I1(frame_65_127_transed_reg[43]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[43]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[43]),
        .O(\stat_rd_data[43]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[43]_i_7 
       (.I0(underrun_error_reg[43]),
        .I1(multicast_frame_transed_reg[43]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[43]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[43]),
        .O(\stat_rd_data[43]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[44]_i_1 
       (.I0(\stat_rd_data[44]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[44]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[44]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_10 
       (.I0(tagged_frame_transed_reg[44]),
        .I1(frame_1024_max_transed_reg[44]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[44]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[44]),
        .O(\stat_rd_data[44]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_11 
       (.I0(multicast_received_good_reg[44]),
        .I1(broadcast_received_good_reg[44]),
        .I2(out[1]),
        .I3(fcs_error_reg[44]),
        .I4(out[0]),
        .I5(frame_received_good_reg[44]),
        .O(\stat_rd_data[44]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_12 
       (.I0(frame_256_511_good_reg[44]),
        .I1(frame_128_255_good_reg[44]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[44]),
        .I4(out[0]),
        .I5(frame_64_good_reg[44]),
        .O(\stat_rd_data[44]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_13 
       (.I0(lt_out_range_reg[44]),
        .I1(control_frame_good_reg[44]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[44]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[44]),
        .O(\stat_rd_data[44]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_14 
       (.I0(oversize_frame_good_reg[44]),
        .I1(unsupported_control_frame_reg[44]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[44]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[44]),
        .O(\stat_rd_data[44]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_2 
       (.I0(\stat_rd_data_reg[44]_i_4_n_0 ),
        .I1(\stat_rd_data[44]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[44]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[44]_i_7_n_0 ),
        .O(\stat_rd_data[44]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_3 
       (.I0(total_bytes_transed_reg[44]),
        .I1(total_bytes_recved_reg[44]),
        .I2(out[1]),
        .I3(fragment_frame_reg[44]),
        .I4(out[0]),
        .I5(undersize_frame_reg[44]),
        .O(\stat_rd_data[44]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[44]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[44]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[44]),
        .I5(pause_frame_transed_reg[44]),
        .O(\stat_rd_data[44]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_6 
       (.I0(frame_128_255_transed_reg[44]),
        .I1(frame_65_127_transed_reg[44]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[44]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[44]),
        .O(\stat_rd_data[44]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[44]_i_7 
       (.I0(underrun_error_reg[44]),
        .I1(multicast_frame_transed_reg[44]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[44]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[44]),
        .O(\stat_rd_data[44]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[45]_i_1 
       (.I0(\stat_rd_data[45]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[45]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[45]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_10 
       (.I0(tagged_frame_transed_reg[45]),
        .I1(frame_1024_max_transed_reg[45]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[45]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[45]),
        .O(\stat_rd_data[45]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_11 
       (.I0(multicast_received_good_reg[45]),
        .I1(broadcast_received_good_reg[45]),
        .I2(out[1]),
        .I3(fcs_error_reg[45]),
        .I4(out[0]),
        .I5(frame_received_good_reg[45]),
        .O(\stat_rd_data[45]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_12 
       (.I0(frame_256_511_good_reg[45]),
        .I1(frame_128_255_good_reg[45]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[45]),
        .I4(out[0]),
        .I5(frame_64_good_reg[45]),
        .O(\stat_rd_data[45]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_13 
       (.I0(lt_out_range_reg[45]),
        .I1(control_frame_good_reg[45]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[45]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[45]),
        .O(\stat_rd_data[45]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_14 
       (.I0(oversize_frame_good_reg[45]),
        .I1(unsupported_control_frame_reg[45]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[45]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[45]),
        .O(\stat_rd_data[45]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_2 
       (.I0(\stat_rd_data_reg[45]_i_4_n_0 ),
        .I1(\stat_rd_data[45]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[45]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[45]_i_7_n_0 ),
        .O(\stat_rd_data[45]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_3 
       (.I0(total_bytes_transed_reg[45]),
        .I1(total_bytes_recved_reg[45]),
        .I2(out[1]),
        .I3(fragment_frame_reg[45]),
        .I4(out[0]),
        .I5(undersize_frame_reg[45]),
        .O(\stat_rd_data[45]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[45]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[45]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[45]),
        .I5(pause_frame_transed_reg[45]),
        .O(\stat_rd_data[45]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_6 
       (.I0(frame_128_255_transed_reg[45]),
        .I1(frame_65_127_transed_reg[45]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[45]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[45]),
        .O(\stat_rd_data[45]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[45]_i_7 
       (.I0(underrun_error_reg[45]),
        .I1(multicast_frame_transed_reg[45]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[45]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[45]),
        .O(\stat_rd_data[45]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[46]_i_1 
       (.I0(\stat_rd_data[46]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[46]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[46]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_10 
       (.I0(tagged_frame_transed_reg[46]),
        .I1(frame_1024_max_transed_reg[46]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[46]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[46]),
        .O(\stat_rd_data[46]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_11 
       (.I0(multicast_received_good_reg[46]),
        .I1(broadcast_received_good_reg[46]),
        .I2(out[1]),
        .I3(fcs_error_reg[46]),
        .I4(out[0]),
        .I5(frame_received_good_reg[46]),
        .O(\stat_rd_data[46]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_12 
       (.I0(frame_256_511_good_reg[46]),
        .I1(frame_128_255_good_reg[46]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[46]),
        .I4(out[0]),
        .I5(frame_64_good_reg[46]),
        .O(\stat_rd_data[46]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_13 
       (.I0(lt_out_range_reg[46]),
        .I1(control_frame_good_reg[46]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[46]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[46]),
        .O(\stat_rd_data[46]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_14 
       (.I0(oversize_frame_good_reg[46]),
        .I1(unsupported_control_frame_reg[46]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[46]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[46]),
        .O(\stat_rd_data[46]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_2 
       (.I0(\stat_rd_data_reg[46]_i_4_n_0 ),
        .I1(\stat_rd_data[46]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[46]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[46]_i_7_n_0 ),
        .O(\stat_rd_data[46]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_3 
       (.I0(total_bytes_transed_reg[46]),
        .I1(total_bytes_recved_reg[46]),
        .I2(out[1]),
        .I3(fragment_frame_reg[46]),
        .I4(out[0]),
        .I5(undersize_frame_reg[46]),
        .O(\stat_rd_data[46]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[46]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[46]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[46]),
        .I5(pause_frame_transed_reg[46]),
        .O(\stat_rd_data[46]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_6 
       (.I0(frame_128_255_transed_reg[46]),
        .I1(frame_65_127_transed_reg[46]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[46]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[46]),
        .O(\stat_rd_data[46]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[46]_i_7 
       (.I0(underrun_error_reg[46]),
        .I1(multicast_frame_transed_reg[46]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[46]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[46]),
        .O(\stat_rd_data[46]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[47]_i_1 
       (.I0(\stat_rd_data[47]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[47]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[47]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_10 
       (.I0(tagged_frame_transed_reg[47]),
        .I1(frame_1024_max_transed_reg[47]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[47]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[47]),
        .O(\stat_rd_data[47]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_11 
       (.I0(multicast_received_good_reg[47]),
        .I1(broadcast_received_good_reg[47]),
        .I2(out[1]),
        .I3(fcs_error_reg[47]),
        .I4(out[0]),
        .I5(frame_received_good_reg[47]),
        .O(\stat_rd_data[47]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_12 
       (.I0(frame_256_511_good_reg[47]),
        .I1(frame_128_255_good_reg[47]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[47]),
        .I4(out[0]),
        .I5(frame_64_good_reg[47]),
        .O(\stat_rd_data[47]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_13 
       (.I0(lt_out_range_reg[47]),
        .I1(control_frame_good_reg[47]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[47]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[47]),
        .O(\stat_rd_data[47]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_14 
       (.I0(oversize_frame_good_reg[47]),
        .I1(unsupported_control_frame_reg[47]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[47]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[47]),
        .O(\stat_rd_data[47]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_2 
       (.I0(\stat_rd_data_reg[47]_i_4_n_0 ),
        .I1(\stat_rd_data[47]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[47]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[47]_i_7_n_0 ),
        .O(\stat_rd_data[47]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_3 
       (.I0(total_bytes_transed_reg[47]),
        .I1(total_bytes_recved_reg[47]),
        .I2(out[1]),
        .I3(fragment_frame_reg[47]),
        .I4(out[0]),
        .I5(undersize_frame_reg[47]),
        .O(\stat_rd_data[47]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[47]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[47]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[47]),
        .I5(pause_frame_transed_reg[47]),
        .O(\stat_rd_data[47]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_6 
       (.I0(frame_128_255_transed_reg[47]),
        .I1(frame_65_127_transed_reg[47]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[47]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[47]),
        .O(\stat_rd_data[47]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[47]_i_7 
       (.I0(underrun_error_reg[47]),
        .I1(multicast_frame_transed_reg[47]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[47]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[47]),
        .O(\stat_rd_data[47]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[48]_i_1 
       (.I0(\stat_rd_data[48]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[48]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[48]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_10 
       (.I0(tagged_frame_transed_reg[48]),
        .I1(frame_1024_max_transed_reg[48]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[48]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[48]),
        .O(\stat_rd_data[48]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_11 
       (.I0(multicast_received_good_reg[48]),
        .I1(broadcast_received_good_reg[48]),
        .I2(out[1]),
        .I3(fcs_error_reg[48]),
        .I4(out[0]),
        .I5(frame_received_good_reg[48]),
        .O(\stat_rd_data[48]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_12 
       (.I0(frame_256_511_good_reg[48]),
        .I1(frame_128_255_good_reg[48]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[48]),
        .I4(out[0]),
        .I5(frame_64_good_reg[48]),
        .O(\stat_rd_data[48]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_13 
       (.I0(lt_out_range_reg[48]),
        .I1(control_frame_good_reg[48]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[48]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[48]),
        .O(\stat_rd_data[48]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_14 
       (.I0(oversize_frame_good_reg[48]),
        .I1(unsupported_control_frame_reg[48]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[48]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[48]),
        .O(\stat_rd_data[48]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_2 
       (.I0(\stat_rd_data_reg[48]_i_4_n_0 ),
        .I1(\stat_rd_data[48]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[48]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[48]_i_7_n_0 ),
        .O(\stat_rd_data[48]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_3 
       (.I0(total_bytes_transed_reg[48]),
        .I1(total_bytes_recved_reg[48]),
        .I2(out[1]),
        .I3(fragment_frame_reg[48]),
        .I4(out[0]),
        .I5(undersize_frame_reg[48]),
        .O(\stat_rd_data[48]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[48]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[48]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[48]),
        .I5(pause_frame_transed_reg[48]),
        .O(\stat_rd_data[48]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_6 
       (.I0(frame_128_255_transed_reg[48]),
        .I1(frame_65_127_transed_reg[48]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[48]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[48]),
        .O(\stat_rd_data[48]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[48]_i_7 
       (.I0(underrun_error_reg[48]),
        .I1(multicast_frame_transed_reg[48]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[48]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[48]),
        .O(\stat_rd_data[48]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[49]_i_1 
       (.I0(\stat_rd_data[49]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[49]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[49]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_10 
       (.I0(tagged_frame_transed_reg[49]),
        .I1(frame_1024_max_transed_reg[49]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[49]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[49]),
        .O(\stat_rd_data[49]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_11 
       (.I0(multicast_received_good_reg[49]),
        .I1(broadcast_received_good_reg[49]),
        .I2(out[1]),
        .I3(fcs_error_reg[49]),
        .I4(out[0]),
        .I5(frame_received_good_reg[49]),
        .O(\stat_rd_data[49]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_12 
       (.I0(frame_256_511_good_reg[49]),
        .I1(frame_128_255_good_reg[49]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[49]),
        .I4(out[0]),
        .I5(frame_64_good_reg[49]),
        .O(\stat_rd_data[49]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_13 
       (.I0(lt_out_range_reg[49]),
        .I1(control_frame_good_reg[49]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[49]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[49]),
        .O(\stat_rd_data[49]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_14 
       (.I0(oversize_frame_good_reg[49]),
        .I1(unsupported_control_frame_reg[49]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[49]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[49]),
        .O(\stat_rd_data[49]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_2 
       (.I0(\stat_rd_data_reg[49]_i_4_n_0 ),
        .I1(\stat_rd_data[49]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[49]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[49]_i_7_n_0 ),
        .O(\stat_rd_data[49]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_3 
       (.I0(total_bytes_transed_reg[49]),
        .I1(total_bytes_recved_reg[49]),
        .I2(out[1]),
        .I3(fragment_frame_reg[49]),
        .I4(out[0]),
        .I5(undersize_frame_reg[49]),
        .O(\stat_rd_data[49]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[49]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[49]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[49]),
        .I5(pause_frame_transed_reg[49]),
        .O(\stat_rd_data[49]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_6 
       (.I0(frame_128_255_transed_reg[49]),
        .I1(frame_65_127_transed_reg[49]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[49]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[49]),
        .O(\stat_rd_data[49]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[49]_i_7 
       (.I0(underrun_error_reg[49]),
        .I1(multicast_frame_transed_reg[49]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[49]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[49]),
        .O(\stat_rd_data[49]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[4]_i_1 
       (.I0(\stat_rd_data[4]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[4]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_10 
       (.I0(tagged_frame_transed_reg[4]),
        .I1(frame_1024_max_transed_reg[4]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[4]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[4]),
        .O(\stat_rd_data[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_11 
       (.I0(multicast_received_good_reg[4]),
        .I1(broadcast_received_good_reg[4]),
        .I2(out[1]),
        .I3(fcs_error_reg[4]),
        .I4(out[0]),
        .I5(frame_received_good_reg[4]),
        .O(\stat_rd_data[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_12 
       (.I0(frame_256_511_good_reg[4]),
        .I1(frame_128_255_good_reg[4]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[4]),
        .I4(out[0]),
        .I5(frame_64_good_reg[4]),
        .O(\stat_rd_data[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_13 
       (.I0(lt_out_range_reg[4]),
        .I1(control_frame_good_reg[4]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[4]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[4]),
        .O(\stat_rd_data[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_14 
       (.I0(oversize_frame_good_reg[4]),
        .I1(unsupported_control_frame_reg[4]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[4]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[4]),
        .O(\stat_rd_data[4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_2 
       (.I0(\stat_rd_data_reg[4]_i_4_n_0 ),
        .I1(\stat_rd_data[4]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[4]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[4]_i_7_n_0 ),
        .O(\stat_rd_data[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_3 
       (.I0(total_bytes_transed_reg[4]),
        .I1(total_bytes_recved_reg[4]),
        .I2(out[1]),
        .I3(fragment_frame_reg[4]),
        .I4(out[0]),
        .I5(undersize_frame_reg[4]),
        .O(\stat_rd_data[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[4]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[4]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[4]),
        .I5(pause_frame_transed_reg[4]),
        .O(\stat_rd_data[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_6 
       (.I0(frame_128_255_transed_reg[4]),
        .I1(frame_65_127_transed_reg[4]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[4]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[4]),
        .O(\stat_rd_data[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[4]_i_7 
       (.I0(underrun_error_reg[4]),
        .I1(multicast_frame_transed_reg[4]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[4]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[4]),
        .O(\stat_rd_data[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[50]_i_1 
       (.I0(\stat_rd_data[50]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[50]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[50]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_10 
       (.I0(tagged_frame_transed_reg[50]),
        .I1(frame_1024_max_transed_reg[50]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[50]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[50]),
        .O(\stat_rd_data[50]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_11 
       (.I0(multicast_received_good_reg[50]),
        .I1(broadcast_received_good_reg[50]),
        .I2(out[1]),
        .I3(fcs_error_reg[50]),
        .I4(out[0]),
        .I5(frame_received_good_reg[50]),
        .O(\stat_rd_data[50]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_12 
       (.I0(frame_256_511_good_reg[50]),
        .I1(frame_128_255_good_reg[50]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[50]),
        .I4(out[0]),
        .I5(frame_64_good_reg[50]),
        .O(\stat_rd_data[50]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_13 
       (.I0(lt_out_range_reg[50]),
        .I1(control_frame_good_reg[50]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[50]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[50]),
        .O(\stat_rd_data[50]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_14 
       (.I0(oversize_frame_good_reg[50]),
        .I1(unsupported_control_frame_reg[50]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[50]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[50]),
        .O(\stat_rd_data[50]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_2 
       (.I0(\stat_rd_data_reg[50]_i_4_n_0 ),
        .I1(\stat_rd_data[50]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[50]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[50]_i_7_n_0 ),
        .O(\stat_rd_data[50]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_3 
       (.I0(total_bytes_transed_reg[50]),
        .I1(total_bytes_recved_reg[50]),
        .I2(out[1]),
        .I3(fragment_frame_reg[50]),
        .I4(out[0]),
        .I5(undersize_frame_reg[50]),
        .O(\stat_rd_data[50]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[50]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[50]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[50]),
        .I5(pause_frame_transed_reg[50]),
        .O(\stat_rd_data[50]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_6 
       (.I0(frame_128_255_transed_reg[50]),
        .I1(frame_65_127_transed_reg[50]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[50]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[50]),
        .O(\stat_rd_data[50]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[50]_i_7 
       (.I0(underrun_error_reg[50]),
        .I1(multicast_frame_transed_reg[50]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[50]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[50]),
        .O(\stat_rd_data[50]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[51]_i_1 
       (.I0(\stat_rd_data[51]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[51]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[51]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_10 
       (.I0(tagged_frame_transed_reg[51]),
        .I1(frame_1024_max_transed_reg[51]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[51]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[51]),
        .O(\stat_rd_data[51]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_11 
       (.I0(multicast_received_good_reg[51]),
        .I1(broadcast_received_good_reg[51]),
        .I2(out[1]),
        .I3(fcs_error_reg[51]),
        .I4(out[0]),
        .I5(frame_received_good_reg[51]),
        .O(\stat_rd_data[51]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_12 
       (.I0(frame_256_511_good_reg[51]),
        .I1(frame_128_255_good_reg[51]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[51]),
        .I4(out[0]),
        .I5(frame_64_good_reg[51]),
        .O(\stat_rd_data[51]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_13 
       (.I0(lt_out_range_reg[51]),
        .I1(control_frame_good_reg[51]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[51]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[51]),
        .O(\stat_rd_data[51]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_14 
       (.I0(oversize_frame_good_reg[51]),
        .I1(unsupported_control_frame_reg[51]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[51]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[51]),
        .O(\stat_rd_data[51]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_2 
       (.I0(\stat_rd_data_reg[51]_i_4_n_0 ),
        .I1(\stat_rd_data[51]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[51]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[51]_i_7_n_0 ),
        .O(\stat_rd_data[51]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_3 
       (.I0(total_bytes_transed_reg[51]),
        .I1(total_bytes_recved_reg[51]),
        .I2(out[1]),
        .I3(fragment_frame_reg[51]),
        .I4(out[0]),
        .I5(undersize_frame_reg[51]),
        .O(\stat_rd_data[51]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[51]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[51]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[51]),
        .I5(pause_frame_transed_reg[51]),
        .O(\stat_rd_data[51]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_6 
       (.I0(frame_128_255_transed_reg[51]),
        .I1(frame_65_127_transed_reg[51]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[51]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[51]),
        .O(\stat_rd_data[51]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[51]_i_7 
       (.I0(underrun_error_reg[51]),
        .I1(multicast_frame_transed_reg[51]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[51]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[51]),
        .O(\stat_rd_data[51]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[52]_i_1 
       (.I0(\stat_rd_data[52]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[52]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[52]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_10 
       (.I0(tagged_frame_transed_reg[52]),
        .I1(frame_1024_max_transed_reg[52]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[52]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[52]),
        .O(\stat_rd_data[52]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_11 
       (.I0(multicast_received_good_reg[52]),
        .I1(broadcast_received_good_reg[52]),
        .I2(out[1]),
        .I3(fcs_error_reg[52]),
        .I4(out[0]),
        .I5(frame_received_good_reg[52]),
        .O(\stat_rd_data[52]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_12 
       (.I0(frame_256_511_good_reg[52]),
        .I1(frame_128_255_good_reg[52]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[52]),
        .I4(out[0]),
        .I5(frame_64_good_reg[52]),
        .O(\stat_rd_data[52]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_13 
       (.I0(lt_out_range_reg[52]),
        .I1(control_frame_good_reg[52]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[52]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[52]),
        .O(\stat_rd_data[52]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_14 
       (.I0(oversize_frame_good_reg[52]),
        .I1(unsupported_control_frame_reg[52]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[52]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[52]),
        .O(\stat_rd_data[52]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_2 
       (.I0(\stat_rd_data_reg[52]_i_4_n_0 ),
        .I1(\stat_rd_data[52]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[52]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[52]_i_7_n_0 ),
        .O(\stat_rd_data[52]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_3 
       (.I0(total_bytes_transed_reg[52]),
        .I1(total_bytes_recved_reg[52]),
        .I2(out[1]),
        .I3(fragment_frame_reg[52]),
        .I4(out[0]),
        .I5(undersize_frame_reg[52]),
        .O(\stat_rd_data[52]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[52]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[52]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[52]),
        .I5(pause_frame_transed_reg[52]),
        .O(\stat_rd_data[52]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_6 
       (.I0(frame_128_255_transed_reg[52]),
        .I1(frame_65_127_transed_reg[52]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[52]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[52]),
        .O(\stat_rd_data[52]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[52]_i_7 
       (.I0(underrun_error_reg[52]),
        .I1(multicast_frame_transed_reg[52]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[52]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[52]),
        .O(\stat_rd_data[52]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[53]_i_1 
       (.I0(\stat_rd_data[53]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[53]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[53]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_10 
       (.I0(tagged_frame_transed_reg[53]),
        .I1(frame_1024_max_transed_reg[53]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[53]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[53]),
        .O(\stat_rd_data[53]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_11 
       (.I0(multicast_received_good_reg[53]),
        .I1(broadcast_received_good_reg[53]),
        .I2(out[1]),
        .I3(fcs_error_reg[53]),
        .I4(out[0]),
        .I5(frame_received_good_reg[53]),
        .O(\stat_rd_data[53]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_12 
       (.I0(frame_256_511_good_reg[53]),
        .I1(frame_128_255_good_reg[53]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[53]),
        .I4(out[0]),
        .I5(frame_64_good_reg[53]),
        .O(\stat_rd_data[53]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_13 
       (.I0(lt_out_range_reg[53]),
        .I1(control_frame_good_reg[53]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[53]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[53]),
        .O(\stat_rd_data[53]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_14 
       (.I0(oversize_frame_good_reg[53]),
        .I1(unsupported_control_frame_reg[53]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[53]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[53]),
        .O(\stat_rd_data[53]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_2 
       (.I0(\stat_rd_data_reg[53]_i_4_n_0 ),
        .I1(\stat_rd_data[53]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[53]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[53]_i_7_n_0 ),
        .O(\stat_rd_data[53]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_3 
       (.I0(total_bytes_transed_reg[53]),
        .I1(total_bytes_recved_reg[53]),
        .I2(out[1]),
        .I3(fragment_frame_reg[53]),
        .I4(out[0]),
        .I5(undersize_frame_reg[53]),
        .O(\stat_rd_data[53]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[53]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[53]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[53]),
        .I5(pause_frame_transed_reg[53]),
        .O(\stat_rd_data[53]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_6 
       (.I0(frame_128_255_transed_reg[53]),
        .I1(frame_65_127_transed_reg[53]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[53]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[53]),
        .O(\stat_rd_data[53]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[53]_i_7 
       (.I0(underrun_error_reg[53]),
        .I1(multicast_frame_transed_reg[53]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[53]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[53]),
        .O(\stat_rd_data[53]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[54]_i_1 
       (.I0(\stat_rd_data[54]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[54]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[54]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_10 
       (.I0(tagged_frame_transed_reg[54]),
        .I1(frame_1024_max_transed_reg[54]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[54]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[54]),
        .O(\stat_rd_data[54]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_11 
       (.I0(multicast_received_good_reg[54]),
        .I1(broadcast_received_good_reg[54]),
        .I2(out[1]),
        .I3(fcs_error_reg[54]),
        .I4(out[0]),
        .I5(frame_received_good_reg[54]),
        .O(\stat_rd_data[54]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_12 
       (.I0(frame_256_511_good_reg[54]),
        .I1(frame_128_255_good_reg[54]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[54]),
        .I4(out[0]),
        .I5(frame_64_good_reg[54]),
        .O(\stat_rd_data[54]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_13 
       (.I0(lt_out_range_reg[54]),
        .I1(control_frame_good_reg[54]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[54]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[54]),
        .O(\stat_rd_data[54]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_14 
       (.I0(oversize_frame_good_reg[54]),
        .I1(unsupported_control_frame_reg[54]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[54]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[54]),
        .O(\stat_rd_data[54]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_2 
       (.I0(\stat_rd_data_reg[54]_i_4_n_0 ),
        .I1(\stat_rd_data[54]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[54]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[54]_i_7_n_0 ),
        .O(\stat_rd_data[54]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_3 
       (.I0(total_bytes_transed_reg[54]),
        .I1(total_bytes_recved_reg[54]),
        .I2(out[1]),
        .I3(fragment_frame_reg[54]),
        .I4(out[0]),
        .I5(undersize_frame_reg[54]),
        .O(\stat_rd_data[54]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[54]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[54]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[54]),
        .I5(pause_frame_transed_reg[54]),
        .O(\stat_rd_data[54]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_6 
       (.I0(frame_128_255_transed_reg[54]),
        .I1(frame_65_127_transed_reg[54]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[54]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[54]),
        .O(\stat_rd_data[54]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[54]_i_7 
       (.I0(underrun_error_reg[54]),
        .I1(multicast_frame_transed_reg[54]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[54]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[54]),
        .O(\stat_rd_data[54]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[55]_i_1 
       (.I0(\stat_rd_data[55]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[55]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[55]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_10 
       (.I0(tagged_frame_transed_reg[55]),
        .I1(frame_1024_max_transed_reg[55]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[55]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[55]),
        .O(\stat_rd_data[55]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_11 
       (.I0(multicast_received_good_reg[55]),
        .I1(broadcast_received_good_reg[55]),
        .I2(out[1]),
        .I3(fcs_error_reg[55]),
        .I4(out[0]),
        .I5(frame_received_good_reg[55]),
        .O(\stat_rd_data[55]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_12 
       (.I0(frame_256_511_good_reg[55]),
        .I1(frame_128_255_good_reg[55]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[55]),
        .I4(out[0]),
        .I5(frame_64_good_reg[55]),
        .O(\stat_rd_data[55]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_13 
       (.I0(lt_out_range_reg[55]),
        .I1(control_frame_good_reg[55]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[55]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[55]),
        .O(\stat_rd_data[55]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_14 
       (.I0(oversize_frame_good_reg[55]),
        .I1(unsupported_control_frame_reg[55]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[55]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[55]),
        .O(\stat_rd_data[55]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_2 
       (.I0(\stat_rd_data_reg[55]_i_4_n_0 ),
        .I1(\stat_rd_data[55]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[55]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[55]_i_7_n_0 ),
        .O(\stat_rd_data[55]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_3 
       (.I0(total_bytes_transed_reg[55]),
        .I1(total_bytes_recved_reg[55]),
        .I2(out[1]),
        .I3(fragment_frame_reg[55]),
        .I4(out[0]),
        .I5(undersize_frame_reg[55]),
        .O(\stat_rd_data[55]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[55]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[55]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[55]),
        .I5(pause_frame_transed_reg[55]),
        .O(\stat_rd_data[55]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_6 
       (.I0(frame_128_255_transed_reg[55]),
        .I1(frame_65_127_transed_reg[55]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[55]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[55]),
        .O(\stat_rd_data[55]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[55]_i_7 
       (.I0(underrun_error_reg[55]),
        .I1(multicast_frame_transed_reg[55]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[55]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[55]),
        .O(\stat_rd_data[55]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[56]_i_1 
       (.I0(\stat_rd_data[56]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[56]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[56]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_10 
       (.I0(tagged_frame_transed_reg[56]),
        .I1(frame_1024_max_transed_reg[56]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[56]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[56]),
        .O(\stat_rd_data[56]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_11 
       (.I0(multicast_received_good_reg[56]),
        .I1(broadcast_received_good_reg[56]),
        .I2(out[1]),
        .I3(fcs_error_reg[56]),
        .I4(out[0]),
        .I5(frame_received_good_reg[56]),
        .O(\stat_rd_data[56]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_12 
       (.I0(frame_256_511_good_reg[56]),
        .I1(frame_128_255_good_reg[56]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[56]),
        .I4(out[0]),
        .I5(frame_64_good_reg[56]),
        .O(\stat_rd_data[56]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_13 
       (.I0(lt_out_range_reg[56]),
        .I1(control_frame_good_reg[56]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[56]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[56]),
        .O(\stat_rd_data[56]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_14 
       (.I0(oversize_frame_good_reg[56]),
        .I1(unsupported_control_frame_reg[56]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[56]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[56]),
        .O(\stat_rd_data[56]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_2 
       (.I0(\stat_rd_data_reg[56]_i_4_n_0 ),
        .I1(\stat_rd_data[56]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[56]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[56]_i_7_n_0 ),
        .O(\stat_rd_data[56]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_3 
       (.I0(total_bytes_transed_reg[56]),
        .I1(total_bytes_recved_reg[56]),
        .I2(out[1]),
        .I3(fragment_frame_reg[56]),
        .I4(out[0]),
        .I5(undersize_frame_reg[56]),
        .O(\stat_rd_data[56]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[56]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[56]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[56]),
        .I5(pause_frame_transed_reg[56]),
        .O(\stat_rd_data[56]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_6 
       (.I0(frame_128_255_transed_reg[56]),
        .I1(frame_65_127_transed_reg[56]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[56]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[56]),
        .O(\stat_rd_data[56]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[56]_i_7 
       (.I0(underrun_error_reg[56]),
        .I1(multicast_frame_transed_reg[56]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[56]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[56]),
        .O(\stat_rd_data[56]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[57]_i_1 
       (.I0(\stat_rd_data[57]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[57]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[57]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_10 
       (.I0(tagged_frame_transed_reg[57]),
        .I1(frame_1024_max_transed_reg[57]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[57]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[57]),
        .O(\stat_rd_data[57]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_11 
       (.I0(multicast_received_good_reg[57]),
        .I1(broadcast_received_good_reg[57]),
        .I2(out[1]),
        .I3(fcs_error_reg[57]),
        .I4(out[0]),
        .I5(frame_received_good_reg[57]),
        .O(\stat_rd_data[57]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_12 
       (.I0(frame_256_511_good_reg[57]),
        .I1(frame_128_255_good_reg[57]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[57]),
        .I4(out[0]),
        .I5(frame_64_good_reg[57]),
        .O(\stat_rd_data[57]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_13 
       (.I0(lt_out_range_reg[57]),
        .I1(control_frame_good_reg[57]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[57]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[57]),
        .O(\stat_rd_data[57]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_14 
       (.I0(oversize_frame_good_reg[57]),
        .I1(unsupported_control_frame_reg[57]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[57]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[57]),
        .O(\stat_rd_data[57]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_2 
       (.I0(\stat_rd_data_reg[57]_i_4_n_0 ),
        .I1(\stat_rd_data[57]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[57]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[57]_i_7_n_0 ),
        .O(\stat_rd_data[57]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_3 
       (.I0(total_bytes_transed_reg[57]),
        .I1(total_bytes_recved_reg[57]),
        .I2(out[1]),
        .I3(fragment_frame_reg[57]),
        .I4(out[0]),
        .I5(undersize_frame_reg[57]),
        .O(\stat_rd_data[57]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[57]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[57]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[57]),
        .I5(pause_frame_transed_reg[57]),
        .O(\stat_rd_data[57]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_6 
       (.I0(frame_128_255_transed_reg[57]),
        .I1(frame_65_127_transed_reg[57]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[57]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[57]),
        .O(\stat_rd_data[57]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[57]_i_7 
       (.I0(underrun_error_reg[57]),
        .I1(multicast_frame_transed_reg[57]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[57]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[57]),
        .O(\stat_rd_data[57]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[58]_i_1 
       (.I0(\stat_rd_data[58]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[58]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[58]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_10 
       (.I0(tagged_frame_transed_reg[58]),
        .I1(frame_1024_max_transed_reg[58]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[58]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[58]),
        .O(\stat_rd_data[58]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_11 
       (.I0(multicast_received_good_reg[58]),
        .I1(broadcast_received_good_reg[58]),
        .I2(out[1]),
        .I3(fcs_error_reg[58]),
        .I4(out[0]),
        .I5(frame_received_good_reg[58]),
        .O(\stat_rd_data[58]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_12 
       (.I0(frame_256_511_good_reg[58]),
        .I1(frame_128_255_good_reg[58]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[58]),
        .I4(out[0]),
        .I5(frame_64_good_reg[58]),
        .O(\stat_rd_data[58]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_13 
       (.I0(lt_out_range_reg[58]),
        .I1(control_frame_good_reg[58]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[58]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[58]),
        .O(\stat_rd_data[58]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_14 
       (.I0(oversize_frame_good_reg[58]),
        .I1(unsupported_control_frame_reg[58]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[58]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[58]),
        .O(\stat_rd_data[58]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_2 
       (.I0(\stat_rd_data_reg[58]_i_4_n_0 ),
        .I1(\stat_rd_data[58]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[58]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[58]_i_7_n_0 ),
        .O(\stat_rd_data[58]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_3 
       (.I0(total_bytes_transed_reg[58]),
        .I1(total_bytes_recved_reg[58]),
        .I2(out[1]),
        .I3(fragment_frame_reg[58]),
        .I4(out[0]),
        .I5(undersize_frame_reg[58]),
        .O(\stat_rd_data[58]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[58]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[58]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[58]),
        .I5(pause_frame_transed_reg[58]),
        .O(\stat_rd_data[58]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_6 
       (.I0(frame_128_255_transed_reg[58]),
        .I1(frame_65_127_transed_reg[58]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[58]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[58]),
        .O(\stat_rd_data[58]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[58]_i_7 
       (.I0(underrun_error_reg[58]),
        .I1(multicast_frame_transed_reg[58]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[58]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[58]),
        .O(\stat_rd_data[58]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[59]_i_1 
       (.I0(\stat_rd_data[59]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[59]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[59]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_10 
       (.I0(tagged_frame_transed_reg[59]),
        .I1(frame_1024_max_transed_reg[59]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[59]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[59]),
        .O(\stat_rd_data[59]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_11 
       (.I0(multicast_received_good_reg[59]),
        .I1(broadcast_received_good_reg[59]),
        .I2(out[1]),
        .I3(fcs_error_reg[59]),
        .I4(out[0]),
        .I5(frame_received_good_reg[59]),
        .O(\stat_rd_data[59]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_12 
       (.I0(frame_256_511_good_reg[59]),
        .I1(frame_128_255_good_reg[59]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[59]),
        .I4(out[0]),
        .I5(frame_64_good_reg[59]),
        .O(\stat_rd_data[59]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_13 
       (.I0(lt_out_range_reg[59]),
        .I1(control_frame_good_reg[59]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[59]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[59]),
        .O(\stat_rd_data[59]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_14 
       (.I0(oversize_frame_good_reg[59]),
        .I1(unsupported_control_frame_reg[59]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[59]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[59]),
        .O(\stat_rd_data[59]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_2 
       (.I0(\stat_rd_data_reg[59]_i_4_n_0 ),
        .I1(\stat_rd_data[59]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[59]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[59]_i_7_n_0 ),
        .O(\stat_rd_data[59]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_3 
       (.I0(total_bytes_transed_reg[59]),
        .I1(total_bytes_recved_reg[59]),
        .I2(out[1]),
        .I3(fragment_frame_reg[59]),
        .I4(out[0]),
        .I5(undersize_frame_reg[59]),
        .O(\stat_rd_data[59]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[59]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[59]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[59]),
        .I5(pause_frame_transed_reg[59]),
        .O(\stat_rd_data[59]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_6 
       (.I0(frame_128_255_transed_reg[59]),
        .I1(frame_65_127_transed_reg[59]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[59]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[59]),
        .O(\stat_rd_data[59]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[59]_i_7 
       (.I0(underrun_error_reg[59]),
        .I1(multicast_frame_transed_reg[59]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[59]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[59]),
        .O(\stat_rd_data[59]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[5]_i_1 
       (.I0(\stat_rd_data[5]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[5]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_10 
       (.I0(tagged_frame_transed_reg[5]),
        .I1(frame_1024_max_transed_reg[5]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[5]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[5]),
        .O(\stat_rd_data[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_11 
       (.I0(multicast_received_good_reg[5]),
        .I1(broadcast_received_good_reg[5]),
        .I2(out[1]),
        .I3(fcs_error_reg[5]),
        .I4(out[0]),
        .I5(frame_received_good_reg[5]),
        .O(\stat_rd_data[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_12 
       (.I0(frame_256_511_good_reg[5]),
        .I1(frame_128_255_good_reg[5]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[5]),
        .I4(out[0]),
        .I5(frame_64_good_reg[5]),
        .O(\stat_rd_data[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_13 
       (.I0(lt_out_range_reg[5]),
        .I1(control_frame_good_reg[5]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[5]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[5]),
        .O(\stat_rd_data[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_14 
       (.I0(oversize_frame_good_reg[5]),
        .I1(unsupported_control_frame_reg[5]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[5]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[5]),
        .O(\stat_rd_data[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_2 
       (.I0(\stat_rd_data_reg[5]_i_4_n_0 ),
        .I1(\stat_rd_data[5]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[5]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[5]_i_7_n_0 ),
        .O(\stat_rd_data[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_3 
       (.I0(total_bytes_transed_reg[5]),
        .I1(total_bytes_recved_reg[5]),
        .I2(out[1]),
        .I3(fragment_frame_reg[5]),
        .I4(out[0]),
        .I5(undersize_frame_reg[5]),
        .O(\stat_rd_data[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[5]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[5]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[5]),
        .I5(pause_frame_transed_reg[5]),
        .O(\stat_rd_data[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_6 
       (.I0(frame_128_255_transed_reg[5]),
        .I1(frame_65_127_transed_reg[5]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[5]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[5]),
        .O(\stat_rd_data[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[5]_i_7 
       (.I0(underrun_error_reg[5]),
        .I1(multicast_frame_transed_reg[5]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[5]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[5]),
        .O(\stat_rd_data[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[60]_i_1 
       (.I0(\stat_rd_data[60]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[60]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[60]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_10 
       (.I0(tagged_frame_transed_reg[60]),
        .I1(frame_1024_max_transed_reg[60]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[60]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[60]),
        .O(\stat_rd_data[60]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_11 
       (.I0(multicast_received_good_reg[60]),
        .I1(broadcast_received_good_reg[60]),
        .I2(out[1]),
        .I3(fcs_error_reg[60]),
        .I4(out[0]),
        .I5(frame_received_good_reg[60]),
        .O(\stat_rd_data[60]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_12 
       (.I0(frame_256_511_good_reg[60]),
        .I1(frame_128_255_good_reg[60]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[60]),
        .I4(out[0]),
        .I5(frame_64_good_reg[60]),
        .O(\stat_rd_data[60]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_13 
       (.I0(lt_out_range_reg[60]),
        .I1(control_frame_good_reg[60]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[60]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[60]),
        .O(\stat_rd_data[60]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_14 
       (.I0(oversize_frame_good_reg[60]),
        .I1(unsupported_control_frame_reg[60]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[60]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[60]),
        .O(\stat_rd_data[60]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_2 
       (.I0(\stat_rd_data_reg[60]_i_4_n_0 ),
        .I1(\stat_rd_data[60]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[60]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[60]_i_7_n_0 ),
        .O(\stat_rd_data[60]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_3 
       (.I0(total_bytes_transed_reg[60]),
        .I1(total_bytes_recved_reg[60]),
        .I2(out[1]),
        .I3(fragment_frame_reg[60]),
        .I4(out[0]),
        .I5(undersize_frame_reg[60]),
        .O(\stat_rd_data[60]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[60]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[60]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[60]),
        .I5(pause_frame_transed_reg[60]),
        .O(\stat_rd_data[60]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_6 
       (.I0(frame_128_255_transed_reg[60]),
        .I1(frame_65_127_transed_reg[60]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[60]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[60]),
        .O(\stat_rd_data[60]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[60]_i_7 
       (.I0(underrun_error_reg[60]),
        .I1(multicast_frame_transed_reg[60]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[60]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[60]),
        .O(\stat_rd_data[60]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[61]_i_1 
       (.I0(\stat_rd_data[61]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[61]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[61]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_10 
       (.I0(tagged_frame_transed_reg[61]),
        .I1(frame_1024_max_transed_reg[61]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[61]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[61]),
        .O(\stat_rd_data[61]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_11 
       (.I0(multicast_received_good_reg[61]),
        .I1(broadcast_received_good_reg[61]),
        .I2(out[1]),
        .I3(fcs_error_reg[61]),
        .I4(out[0]),
        .I5(frame_received_good_reg[61]),
        .O(\stat_rd_data[61]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_12 
       (.I0(frame_256_511_good_reg[61]),
        .I1(frame_128_255_good_reg[61]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[61]),
        .I4(out[0]),
        .I5(frame_64_good_reg[61]),
        .O(\stat_rd_data[61]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_13 
       (.I0(lt_out_range_reg[61]),
        .I1(control_frame_good_reg[61]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[61]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[61]),
        .O(\stat_rd_data[61]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_14 
       (.I0(oversize_frame_good_reg[61]),
        .I1(unsupported_control_frame_reg[61]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[61]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[61]),
        .O(\stat_rd_data[61]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_2 
       (.I0(\stat_rd_data_reg[61]_i_4_n_0 ),
        .I1(\stat_rd_data[61]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[61]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[61]_i_7_n_0 ),
        .O(\stat_rd_data[61]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_3 
       (.I0(total_bytes_transed_reg[61]),
        .I1(total_bytes_recved_reg[61]),
        .I2(out[1]),
        .I3(fragment_frame_reg[61]),
        .I4(out[0]),
        .I5(undersize_frame_reg[61]),
        .O(\stat_rd_data[61]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[61]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[61]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[61]),
        .I5(pause_frame_transed_reg[61]),
        .O(\stat_rd_data[61]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_6 
       (.I0(frame_128_255_transed_reg[61]),
        .I1(frame_65_127_transed_reg[61]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[61]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[61]),
        .O(\stat_rd_data[61]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[61]_i_7 
       (.I0(underrun_error_reg[61]),
        .I1(multicast_frame_transed_reg[61]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[61]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[61]),
        .O(\stat_rd_data[61]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[62]_i_1 
       (.I0(\stat_rd_data[62]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[62]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[62]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_10 
       (.I0(tagged_frame_transed_reg[62]),
        .I1(frame_1024_max_transed_reg[62]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[62]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[62]),
        .O(\stat_rd_data[62]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_11 
       (.I0(multicast_received_good_reg[62]),
        .I1(broadcast_received_good_reg[62]),
        .I2(out[1]),
        .I3(fcs_error_reg[62]),
        .I4(out[0]),
        .I5(frame_received_good_reg[62]),
        .O(\stat_rd_data[62]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_12 
       (.I0(frame_256_511_good_reg[62]),
        .I1(frame_128_255_good_reg[62]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[62]),
        .I4(out[0]),
        .I5(frame_64_good_reg[62]),
        .O(\stat_rd_data[62]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_13 
       (.I0(lt_out_range_reg[62]),
        .I1(control_frame_good_reg[62]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[62]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[62]),
        .O(\stat_rd_data[62]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_14 
       (.I0(oversize_frame_good_reg[62]),
        .I1(unsupported_control_frame_reg[62]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[62]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[62]),
        .O(\stat_rd_data[62]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_2 
       (.I0(\stat_rd_data_reg[62]_i_4_n_0 ),
        .I1(\stat_rd_data[62]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[62]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[62]_i_7_n_0 ),
        .O(\stat_rd_data[62]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_3 
       (.I0(total_bytes_transed_reg[62]),
        .I1(total_bytes_recved_reg[62]),
        .I2(out[1]),
        .I3(fragment_frame_reg[62]),
        .I4(out[0]),
        .I5(undersize_frame_reg[62]),
        .O(\stat_rd_data[62]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[62]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[62]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[62]),
        .I5(pause_frame_transed_reg[62]),
        .O(\stat_rd_data[62]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_6 
       (.I0(frame_128_255_transed_reg[62]),
        .I1(frame_65_127_transed_reg[62]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[62]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[62]),
        .O(\stat_rd_data[62]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[62]_i_7 
       (.I0(underrun_error_reg[62]),
        .I1(multicast_frame_transed_reg[62]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[62]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[62]),
        .O(\stat_rd_data[62]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \stat_rd_data[63]_i_1 
       (.I0(out[9]),
        .I1(\stat_rd_data_reg[63]_0 ),
        .I2(\stat_rd_data_reg[63]_1 ),
        .O(\stat_rd_data[63]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat_rd_data[63]_i_10 
       (.I0(out[3]),
        .I1(out[5]),
        .O(\stat_rd_data[63]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_11 
       (.I0(frame_128_255_transed_reg[63]),
        .I1(frame_65_127_transed_reg[63]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[63]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[63]),
        .O(\stat_rd_data[63]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \stat_rd_data[63]_i_12 
       (.I0(out[5]),
        .I1(out[2]),
        .I2(out[3]),
        .O(\stat_rd_data[63]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_13 
       (.I0(underrun_error_reg[63]),
        .I1(multicast_frame_transed_reg[63]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[63]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[63]),
        .O(\stat_rd_data[63]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_16 
       (.I0(tagged_frame_transed_reg[63]),
        .I1(frame_1024_max_transed_reg[63]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[63]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[63]),
        .O(\stat_rd_data[63]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_17 
       (.I0(multicast_received_good_reg[63]),
        .I1(broadcast_received_good_reg[63]),
        .I2(out[1]),
        .I3(fcs_error_reg[63]),
        .I4(out[0]),
        .I5(frame_received_good_reg[63]),
        .O(\stat_rd_data[63]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_18 
       (.I0(frame_256_511_good_reg[63]),
        .I1(frame_128_255_good_reg[63]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[63]),
        .I4(out[0]),
        .I5(frame_64_good_reg[63]),
        .O(\stat_rd_data[63]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_19 
       (.I0(lt_out_range_reg[63]),
        .I1(control_frame_good_reg[63]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[63]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[63]),
        .O(\stat_rd_data[63]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[63]_i_2 
       (.I0(\stat_rd_data[63]_i_3_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[63]_i_5_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[63]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_20 
       (.I0(oversize_frame_good_reg[63]),
        .I1(unsupported_control_frame_reg[63]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[63]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[63]),
        .O(\stat_rd_data[63]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_3 
       (.I0(\stat_rd_data_reg[63]_i_8_n_0 ),
        .I1(\stat_rd_data[63]_i_9_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[63]_i_11_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[63]_i_13_n_0 ),
        .O(\stat_rd_data[63]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat_rd_data[63]_i_4 
       (.I0(out[3]),
        .I1(out[5]),
        .O(\stat_rd_data[63]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[63]_i_5 
       (.I0(total_bytes_transed_reg[63]),
        .I1(total_bytes_recved_reg[63]),
        .I2(out[1]),
        .I3(fragment_frame_reg[63]),
        .I4(out[0]),
        .I5(undersize_frame_reg[63]),
        .O(\stat_rd_data[63]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \stat_rd_data[63]_i_6 
       (.I0(out[5]),
        .I1(out[3]),
        .I2(out[2]),
        .O(\stat_rd_data[63]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat_rd_data[63]_i_7 
       (.I0(out[7]),
        .I1(out[6]),
        .O(\stat_rd_data[63]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[63]_i_9 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[63]_i_16_n_0 ),
        .I4(oversize_frame_transed_reg[63]),
        .I5(pause_frame_transed_reg[63]),
        .O(\stat_rd_data[63]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[6]_i_1 
       (.I0(\stat_rd_data[6]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[6]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_10 
       (.I0(tagged_frame_transed_reg[6]),
        .I1(frame_1024_max_transed_reg[6]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[6]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[6]),
        .O(\stat_rd_data[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_11 
       (.I0(multicast_received_good_reg[6]),
        .I1(broadcast_received_good_reg[6]),
        .I2(out[1]),
        .I3(fcs_error_reg[6]),
        .I4(out[0]),
        .I5(frame_received_good_reg[6]),
        .O(\stat_rd_data[6]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_12 
       (.I0(frame_256_511_good_reg[6]),
        .I1(frame_128_255_good_reg[6]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[6]),
        .I4(out[0]),
        .I5(frame_64_good_reg[6]),
        .O(\stat_rd_data[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_13 
       (.I0(lt_out_range_reg[6]),
        .I1(control_frame_good_reg[6]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[6]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[6]),
        .O(\stat_rd_data[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_14 
       (.I0(oversize_frame_good_reg[6]),
        .I1(unsupported_control_frame_reg[6]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[6]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[6]),
        .O(\stat_rd_data[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_2 
       (.I0(\stat_rd_data_reg[6]_i_4_n_0 ),
        .I1(\stat_rd_data[6]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[6]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[6]_i_7_n_0 ),
        .O(\stat_rd_data[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_3 
       (.I0(total_bytes_transed_reg[6]),
        .I1(total_bytes_recved_reg[6]),
        .I2(out[1]),
        .I3(fragment_frame_reg[6]),
        .I4(out[0]),
        .I5(undersize_frame_reg[6]),
        .O(\stat_rd_data[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[6]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[6]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[6]),
        .I5(pause_frame_transed_reg[6]),
        .O(\stat_rd_data[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_6 
       (.I0(frame_128_255_transed_reg[6]),
        .I1(frame_65_127_transed_reg[6]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[6]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[6]),
        .O(\stat_rd_data[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[6]_i_7 
       (.I0(underrun_error_reg[6]),
        .I1(multicast_frame_transed_reg[6]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[6]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[6]),
        .O(\stat_rd_data[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[7]_i_1 
       (.I0(\stat_rd_data[7]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[7]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_10 
       (.I0(tagged_frame_transed_reg[7]),
        .I1(frame_1024_max_transed_reg[7]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[7]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[7]),
        .O(\stat_rd_data[7]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_11 
       (.I0(multicast_received_good_reg[7]),
        .I1(broadcast_received_good_reg[7]),
        .I2(out[1]),
        .I3(fcs_error_reg[7]),
        .I4(out[0]),
        .I5(frame_received_good_reg[7]),
        .O(\stat_rd_data[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_12 
       (.I0(frame_256_511_good_reg[7]),
        .I1(frame_128_255_good_reg[7]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[7]),
        .I4(out[0]),
        .I5(frame_64_good_reg[7]),
        .O(\stat_rd_data[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_13 
       (.I0(lt_out_range_reg[7]),
        .I1(control_frame_good_reg[7]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[7]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[7]),
        .O(\stat_rd_data[7]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_14 
       (.I0(oversize_frame_good_reg[7]),
        .I1(unsupported_control_frame_reg[7]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[7]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[7]),
        .O(\stat_rd_data[7]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_2 
       (.I0(\stat_rd_data_reg[7]_i_4_n_0 ),
        .I1(\stat_rd_data[7]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[7]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[7]_i_7_n_0 ),
        .O(\stat_rd_data[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_3 
       (.I0(total_bytes_transed_reg[7]),
        .I1(total_bytes_recved_reg[7]),
        .I2(out[1]),
        .I3(fragment_frame_reg[7]),
        .I4(out[0]),
        .I5(undersize_frame_reg[7]),
        .O(\stat_rd_data[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[7]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[7]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[7]),
        .I5(pause_frame_transed_reg[7]),
        .O(\stat_rd_data[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_6 
       (.I0(frame_128_255_transed_reg[7]),
        .I1(frame_65_127_transed_reg[7]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[7]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[7]),
        .O(\stat_rd_data[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[7]_i_7 
       (.I0(underrun_error_reg[7]),
        .I1(multicast_frame_transed_reg[7]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[7]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[7]),
        .O(\stat_rd_data[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[8]_i_1 
       (.I0(\stat_rd_data[8]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[8]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_10 
       (.I0(tagged_frame_transed_reg[8]),
        .I1(frame_1024_max_transed_reg[8]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[8]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[8]),
        .O(\stat_rd_data[8]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_11 
       (.I0(multicast_received_good_reg[8]),
        .I1(broadcast_received_good_reg[8]),
        .I2(out[1]),
        .I3(fcs_error_reg[8]),
        .I4(out[0]),
        .I5(frame_received_good_reg[8]),
        .O(\stat_rd_data[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_12 
       (.I0(frame_256_511_good_reg[8]),
        .I1(frame_128_255_good_reg[8]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[8]),
        .I4(out[0]),
        .I5(frame_64_good_reg[8]),
        .O(\stat_rd_data[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_13 
       (.I0(lt_out_range_reg[8]),
        .I1(control_frame_good_reg[8]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[8]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[8]),
        .O(\stat_rd_data[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_14 
       (.I0(oversize_frame_good_reg[8]),
        .I1(unsupported_control_frame_reg[8]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[8]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[8]),
        .O(\stat_rd_data[8]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_2 
       (.I0(\stat_rd_data_reg[8]_i_4_n_0 ),
        .I1(\stat_rd_data[8]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[8]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[8]_i_7_n_0 ),
        .O(\stat_rd_data[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_3 
       (.I0(total_bytes_transed_reg[8]),
        .I1(total_bytes_recved_reg[8]),
        .I2(out[1]),
        .I3(fragment_frame_reg[8]),
        .I4(out[0]),
        .I5(undersize_frame_reg[8]),
        .O(\stat_rd_data[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[8]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[8]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[8]),
        .I5(pause_frame_transed_reg[8]),
        .O(\stat_rd_data[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_6 
       (.I0(frame_128_255_transed_reg[8]),
        .I1(frame_65_127_transed_reg[8]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[8]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[8]),
        .O(\stat_rd_data[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[8]_i_7 
       (.I0(underrun_error_reg[8]),
        .I1(multicast_frame_transed_reg[8]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[8]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[8]),
        .O(\stat_rd_data[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222E22)) 
    \stat_rd_data[9]_i_1 
       (.I0(\stat_rd_data[9]_i_2_n_0 ),
        .I1(out[4]),
        .I2(\stat_rd_data[63]_i_4_n_0 ),
        .I3(\stat_rd_data[9]_i_3_n_0 ),
        .I4(\stat_rd_data[63]_i_6_n_0 ),
        .I5(\stat_rd_data[63]_i_7_n_0 ),
        .O(p_0_in[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_10 
       (.I0(tagged_frame_transed_reg[9]),
        .I1(frame_1024_max_transed_reg[9]),
        .I2(out[1]),
        .I3(frame_512_1023_transed_reg[9]),
        .I4(out[0]),
        .I5(frame_256_511_transed_reg[9]),
        .O(\stat_rd_data[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_11 
       (.I0(multicast_received_good_reg[9]),
        .I1(broadcast_received_good_reg[9]),
        .I2(out[1]),
        .I3(fcs_error_reg[9]),
        .I4(out[0]),
        .I5(frame_received_good_reg[9]),
        .O(\stat_rd_data[9]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_12 
       (.I0(frame_256_511_good_reg[9]),
        .I1(frame_128_255_good_reg[9]),
        .I2(out[1]),
        .I3(frame_65_127_good_reg[9]),
        .I4(out[0]),
        .I5(frame_64_good_reg[9]),
        .O(\stat_rd_data[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_13 
       (.I0(lt_out_range_reg[9]),
        .I1(control_frame_good_reg[9]),
        .I2(out[1]),
        .I3(frame_1024_max_good_reg[9]),
        .I4(out[0]),
        .I5(frame_512_1023_good_reg[9]),
        .O(\stat_rd_data[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_14 
       (.I0(oversize_frame_good_reg[9]),
        .I1(unsupported_control_frame_reg[9]),
        .I2(out[1]),
        .I3(pause_frame_good_reg[9]),
        .I4(out[0]),
        .I5(tagged_frame_good_reg[9]),
        .O(\stat_rd_data[9]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_2 
       (.I0(\stat_rd_data_reg[9]_i_4_n_0 ),
        .I1(\stat_rd_data[9]_i_5_n_0 ),
        .I2(\stat_rd_data[63]_i_10_n_0 ),
        .I3(\stat_rd_data[9]_i_6_n_0 ),
        .I4(\stat_rd_data[63]_i_12_n_0 ),
        .I5(\stat_rd_data[9]_i_7_n_0 ),
        .O(\stat_rd_data[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_3 
       (.I0(total_bytes_transed_reg[9]),
        .I1(total_bytes_recved_reg[9]),
        .I2(out[1]),
        .I3(fragment_frame_reg[9]),
        .I4(out[0]),
        .I5(undersize_frame_reg[9]),
        .O(\stat_rd_data[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5F0A57025D085500)) 
    \stat_rd_data[9]_i_5 
       (.I0(out[2]),
        .I1(out[0]),
        .I2(out[1]),
        .I3(\stat_rd_data[9]_i_10_n_0 ),
        .I4(oversize_frame_transed_reg[9]),
        .I5(pause_frame_transed_reg[9]),
        .O(\stat_rd_data[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_6 
       (.I0(frame_128_255_transed_reg[9]),
        .I1(frame_65_127_transed_reg[9]),
        .I2(out[1]),
        .I3(frame_64_transed_reg[9]),
        .I4(out[0]),
        .I5(control_frame_transed_reg[9]),
        .O(\stat_rd_data[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \stat_rd_data[9]_i_7 
       (.I0(underrun_error_reg[9]),
        .I1(multicast_frame_transed_reg[9]),
        .I2(out[1]),
        .I3(broadcast_frame_transed_reg[9]),
        .I4(out[0]),
        .I5(good_frame_transed_reg[9]),
        .O(\stat_rd_data[9]_i_7_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[0] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[0]),
        .Q(stat_rd_data[0]));
  MUXF8 \stat_rd_data_reg[0]_i_4 
       (.I0(\stat_rd_data_reg[0]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[0]_i_9_n_0 ),
        .O(\stat_rd_data_reg[0]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[0]_i_8 
       (.I0(\stat_rd_data[0]_i_11_n_0 ),
        .I1(\stat_rd_data[0]_i_12_n_0 ),
        .O(\stat_rd_data_reg[0]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[0]_i_9 
       (.I0(\stat_rd_data[0]_i_13_n_0 ),
        .I1(\stat_rd_data[0]_i_14_n_0 ),
        .O(\stat_rd_data_reg[0]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[10] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[10]),
        .Q(stat_rd_data[10]));
  MUXF8 \stat_rd_data_reg[10]_i_4 
       (.I0(\stat_rd_data_reg[10]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[10]_i_9_n_0 ),
        .O(\stat_rd_data_reg[10]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[10]_i_8 
       (.I0(\stat_rd_data[10]_i_11_n_0 ),
        .I1(\stat_rd_data[10]_i_12_n_0 ),
        .O(\stat_rd_data_reg[10]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[10]_i_9 
       (.I0(\stat_rd_data[10]_i_13_n_0 ),
        .I1(\stat_rd_data[10]_i_14_n_0 ),
        .O(\stat_rd_data_reg[10]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[11] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[11]),
        .Q(stat_rd_data[11]));
  MUXF8 \stat_rd_data_reg[11]_i_4 
       (.I0(\stat_rd_data_reg[11]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[11]_i_9_n_0 ),
        .O(\stat_rd_data_reg[11]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[11]_i_8 
       (.I0(\stat_rd_data[11]_i_11_n_0 ),
        .I1(\stat_rd_data[11]_i_12_n_0 ),
        .O(\stat_rd_data_reg[11]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[11]_i_9 
       (.I0(\stat_rd_data[11]_i_13_n_0 ),
        .I1(\stat_rd_data[11]_i_14_n_0 ),
        .O(\stat_rd_data_reg[11]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[12] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[12]),
        .Q(stat_rd_data[12]));
  MUXF8 \stat_rd_data_reg[12]_i_4 
       (.I0(\stat_rd_data_reg[12]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[12]_i_9_n_0 ),
        .O(\stat_rd_data_reg[12]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[12]_i_8 
       (.I0(\stat_rd_data[12]_i_11_n_0 ),
        .I1(\stat_rd_data[12]_i_12_n_0 ),
        .O(\stat_rd_data_reg[12]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[12]_i_9 
       (.I0(\stat_rd_data[12]_i_13_n_0 ),
        .I1(\stat_rd_data[12]_i_14_n_0 ),
        .O(\stat_rd_data_reg[12]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[13] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[13]),
        .Q(stat_rd_data[13]));
  MUXF8 \stat_rd_data_reg[13]_i_4 
       (.I0(\stat_rd_data_reg[13]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[13]_i_9_n_0 ),
        .O(\stat_rd_data_reg[13]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[13]_i_8 
       (.I0(\stat_rd_data[13]_i_11_n_0 ),
        .I1(\stat_rd_data[13]_i_12_n_0 ),
        .O(\stat_rd_data_reg[13]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[13]_i_9 
       (.I0(\stat_rd_data[13]_i_13_n_0 ),
        .I1(\stat_rd_data[13]_i_14_n_0 ),
        .O(\stat_rd_data_reg[13]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[14] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[14]),
        .Q(stat_rd_data[14]));
  MUXF8 \stat_rd_data_reg[14]_i_4 
       (.I0(\stat_rd_data_reg[14]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[14]_i_9_n_0 ),
        .O(\stat_rd_data_reg[14]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[14]_i_8 
       (.I0(\stat_rd_data[14]_i_11_n_0 ),
        .I1(\stat_rd_data[14]_i_12_n_0 ),
        .O(\stat_rd_data_reg[14]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[14]_i_9 
       (.I0(\stat_rd_data[14]_i_13_n_0 ),
        .I1(\stat_rd_data[14]_i_14_n_0 ),
        .O(\stat_rd_data_reg[14]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[15] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[15]),
        .Q(stat_rd_data[15]));
  MUXF8 \stat_rd_data_reg[15]_i_4 
       (.I0(\stat_rd_data_reg[15]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[15]_i_9_n_0 ),
        .O(\stat_rd_data_reg[15]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[15]_i_8 
       (.I0(\stat_rd_data[15]_i_11_n_0 ),
        .I1(\stat_rd_data[15]_i_12_n_0 ),
        .O(\stat_rd_data_reg[15]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[15]_i_9 
       (.I0(\stat_rd_data[15]_i_13_n_0 ),
        .I1(\stat_rd_data[15]_i_14_n_0 ),
        .O(\stat_rd_data_reg[15]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[16] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[16]),
        .Q(stat_rd_data[16]));
  MUXF8 \stat_rd_data_reg[16]_i_4 
       (.I0(\stat_rd_data_reg[16]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[16]_i_9_n_0 ),
        .O(\stat_rd_data_reg[16]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[16]_i_8 
       (.I0(\stat_rd_data[16]_i_11_n_0 ),
        .I1(\stat_rd_data[16]_i_12_n_0 ),
        .O(\stat_rd_data_reg[16]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[16]_i_9 
       (.I0(\stat_rd_data[16]_i_13_n_0 ),
        .I1(\stat_rd_data[16]_i_14_n_0 ),
        .O(\stat_rd_data_reg[16]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[17] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[17]),
        .Q(stat_rd_data[17]));
  MUXF8 \stat_rd_data_reg[17]_i_4 
       (.I0(\stat_rd_data_reg[17]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[17]_i_9_n_0 ),
        .O(\stat_rd_data_reg[17]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[17]_i_8 
       (.I0(\stat_rd_data[17]_i_11_n_0 ),
        .I1(\stat_rd_data[17]_i_12_n_0 ),
        .O(\stat_rd_data_reg[17]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[17]_i_9 
       (.I0(\stat_rd_data[17]_i_13_n_0 ),
        .I1(\stat_rd_data[17]_i_14_n_0 ),
        .O(\stat_rd_data_reg[17]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[18] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[18]),
        .Q(stat_rd_data[18]));
  MUXF8 \stat_rd_data_reg[18]_i_4 
       (.I0(\stat_rd_data_reg[18]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[18]_i_9_n_0 ),
        .O(\stat_rd_data_reg[18]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[18]_i_8 
       (.I0(\stat_rd_data[18]_i_11_n_0 ),
        .I1(\stat_rd_data[18]_i_12_n_0 ),
        .O(\stat_rd_data_reg[18]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[18]_i_9 
       (.I0(\stat_rd_data[18]_i_13_n_0 ),
        .I1(\stat_rd_data[18]_i_14_n_0 ),
        .O(\stat_rd_data_reg[18]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[19] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[19]),
        .Q(stat_rd_data[19]));
  MUXF8 \stat_rd_data_reg[19]_i_4 
       (.I0(\stat_rd_data_reg[19]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[19]_i_9_n_0 ),
        .O(\stat_rd_data_reg[19]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[19]_i_8 
       (.I0(\stat_rd_data[19]_i_11_n_0 ),
        .I1(\stat_rd_data[19]_i_12_n_0 ),
        .O(\stat_rd_data_reg[19]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[19]_i_9 
       (.I0(\stat_rd_data[19]_i_13_n_0 ),
        .I1(\stat_rd_data[19]_i_14_n_0 ),
        .O(\stat_rd_data_reg[19]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[1] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[1]),
        .Q(stat_rd_data[1]));
  MUXF8 \stat_rd_data_reg[1]_i_4 
       (.I0(\stat_rd_data_reg[1]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[1]_i_9_n_0 ),
        .O(\stat_rd_data_reg[1]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[1]_i_8 
       (.I0(\stat_rd_data[1]_i_11_n_0 ),
        .I1(\stat_rd_data[1]_i_12_n_0 ),
        .O(\stat_rd_data_reg[1]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[1]_i_9 
       (.I0(\stat_rd_data[1]_i_13_n_0 ),
        .I1(\stat_rd_data[1]_i_14_n_0 ),
        .O(\stat_rd_data_reg[1]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[20] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[20]),
        .Q(stat_rd_data[20]));
  MUXF8 \stat_rd_data_reg[20]_i_4 
       (.I0(\stat_rd_data_reg[20]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[20]_i_9_n_0 ),
        .O(\stat_rd_data_reg[20]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[20]_i_8 
       (.I0(\stat_rd_data[20]_i_11_n_0 ),
        .I1(\stat_rd_data[20]_i_12_n_0 ),
        .O(\stat_rd_data_reg[20]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[20]_i_9 
       (.I0(\stat_rd_data[20]_i_13_n_0 ),
        .I1(\stat_rd_data[20]_i_14_n_0 ),
        .O(\stat_rd_data_reg[20]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[21] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[21]),
        .Q(stat_rd_data[21]));
  MUXF8 \stat_rd_data_reg[21]_i_4 
       (.I0(\stat_rd_data_reg[21]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[21]_i_9_n_0 ),
        .O(\stat_rd_data_reg[21]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[21]_i_8 
       (.I0(\stat_rd_data[21]_i_11_n_0 ),
        .I1(\stat_rd_data[21]_i_12_n_0 ),
        .O(\stat_rd_data_reg[21]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[21]_i_9 
       (.I0(\stat_rd_data[21]_i_13_n_0 ),
        .I1(\stat_rd_data[21]_i_14_n_0 ),
        .O(\stat_rd_data_reg[21]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[22] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[22]),
        .Q(stat_rd_data[22]));
  MUXF8 \stat_rd_data_reg[22]_i_4 
       (.I0(\stat_rd_data_reg[22]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[22]_i_9_n_0 ),
        .O(\stat_rd_data_reg[22]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[22]_i_8 
       (.I0(\stat_rd_data[22]_i_11_n_0 ),
        .I1(\stat_rd_data[22]_i_12_n_0 ),
        .O(\stat_rd_data_reg[22]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[22]_i_9 
       (.I0(\stat_rd_data[22]_i_13_n_0 ),
        .I1(\stat_rd_data[22]_i_14_n_0 ),
        .O(\stat_rd_data_reg[22]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[23] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[23]),
        .Q(stat_rd_data[23]));
  MUXF8 \stat_rd_data_reg[23]_i_4 
       (.I0(\stat_rd_data_reg[23]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[23]_i_9_n_0 ),
        .O(\stat_rd_data_reg[23]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[23]_i_8 
       (.I0(\stat_rd_data[23]_i_11_n_0 ),
        .I1(\stat_rd_data[23]_i_12_n_0 ),
        .O(\stat_rd_data_reg[23]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[23]_i_9 
       (.I0(\stat_rd_data[23]_i_13_n_0 ),
        .I1(\stat_rd_data[23]_i_14_n_0 ),
        .O(\stat_rd_data_reg[23]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[24] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[24]),
        .Q(stat_rd_data[24]));
  MUXF8 \stat_rd_data_reg[24]_i_4 
       (.I0(\stat_rd_data_reg[24]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[24]_i_9_n_0 ),
        .O(\stat_rd_data_reg[24]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[24]_i_8 
       (.I0(\stat_rd_data[24]_i_11_n_0 ),
        .I1(\stat_rd_data[24]_i_12_n_0 ),
        .O(\stat_rd_data_reg[24]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[24]_i_9 
       (.I0(\stat_rd_data[24]_i_13_n_0 ),
        .I1(\stat_rd_data[24]_i_14_n_0 ),
        .O(\stat_rd_data_reg[24]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[25] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[25]),
        .Q(stat_rd_data[25]));
  MUXF8 \stat_rd_data_reg[25]_i_4 
       (.I0(\stat_rd_data_reg[25]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[25]_i_9_n_0 ),
        .O(\stat_rd_data_reg[25]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[25]_i_8 
       (.I0(\stat_rd_data[25]_i_11_n_0 ),
        .I1(\stat_rd_data[25]_i_12_n_0 ),
        .O(\stat_rd_data_reg[25]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[25]_i_9 
       (.I0(\stat_rd_data[25]_i_13_n_0 ),
        .I1(\stat_rd_data[25]_i_14_n_0 ),
        .O(\stat_rd_data_reg[25]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[26] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[26]),
        .Q(stat_rd_data[26]));
  MUXF8 \stat_rd_data_reg[26]_i_4 
       (.I0(\stat_rd_data_reg[26]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[26]_i_9_n_0 ),
        .O(\stat_rd_data_reg[26]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[26]_i_8 
       (.I0(\stat_rd_data[26]_i_11_n_0 ),
        .I1(\stat_rd_data[26]_i_12_n_0 ),
        .O(\stat_rd_data_reg[26]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[26]_i_9 
       (.I0(\stat_rd_data[26]_i_13_n_0 ),
        .I1(\stat_rd_data[26]_i_14_n_0 ),
        .O(\stat_rd_data_reg[26]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[27] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[27]),
        .Q(stat_rd_data[27]));
  MUXF8 \stat_rd_data_reg[27]_i_4 
       (.I0(\stat_rd_data_reg[27]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[27]_i_9_n_0 ),
        .O(\stat_rd_data_reg[27]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[27]_i_8 
       (.I0(\stat_rd_data[27]_i_11_n_0 ),
        .I1(\stat_rd_data[27]_i_12_n_0 ),
        .O(\stat_rd_data_reg[27]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[27]_i_9 
       (.I0(\stat_rd_data[27]_i_13_n_0 ),
        .I1(\stat_rd_data[27]_i_14_n_0 ),
        .O(\stat_rd_data_reg[27]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[28] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[28]),
        .Q(stat_rd_data[28]));
  MUXF8 \stat_rd_data_reg[28]_i_4 
       (.I0(\stat_rd_data_reg[28]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[28]_i_9_n_0 ),
        .O(\stat_rd_data_reg[28]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[28]_i_8 
       (.I0(\stat_rd_data[28]_i_11_n_0 ),
        .I1(\stat_rd_data[28]_i_12_n_0 ),
        .O(\stat_rd_data_reg[28]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[28]_i_9 
       (.I0(\stat_rd_data[28]_i_13_n_0 ),
        .I1(\stat_rd_data[28]_i_14_n_0 ),
        .O(\stat_rd_data_reg[28]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[29] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[29]),
        .Q(stat_rd_data[29]));
  MUXF8 \stat_rd_data_reg[29]_i_4 
       (.I0(\stat_rd_data_reg[29]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[29]_i_9_n_0 ),
        .O(\stat_rd_data_reg[29]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[29]_i_8 
       (.I0(\stat_rd_data[29]_i_11_n_0 ),
        .I1(\stat_rd_data[29]_i_12_n_0 ),
        .O(\stat_rd_data_reg[29]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[29]_i_9 
       (.I0(\stat_rd_data[29]_i_13_n_0 ),
        .I1(\stat_rd_data[29]_i_14_n_0 ),
        .O(\stat_rd_data_reg[29]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[2] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[2]),
        .Q(stat_rd_data[2]));
  MUXF8 \stat_rd_data_reg[2]_i_4 
       (.I0(\stat_rd_data_reg[2]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[2]_i_9_n_0 ),
        .O(\stat_rd_data_reg[2]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[2]_i_8 
       (.I0(\stat_rd_data[2]_i_11_n_0 ),
        .I1(\stat_rd_data[2]_i_12_n_0 ),
        .O(\stat_rd_data_reg[2]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[2]_i_9 
       (.I0(\stat_rd_data[2]_i_13_n_0 ),
        .I1(\stat_rd_data[2]_i_14_n_0 ),
        .O(\stat_rd_data_reg[2]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[30] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[30]),
        .Q(stat_rd_data[30]));
  MUXF8 \stat_rd_data_reg[30]_i_4 
       (.I0(\stat_rd_data_reg[30]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[30]_i_9_n_0 ),
        .O(\stat_rd_data_reg[30]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[30]_i_8 
       (.I0(\stat_rd_data[30]_i_11_n_0 ),
        .I1(\stat_rd_data[30]_i_12_n_0 ),
        .O(\stat_rd_data_reg[30]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[30]_i_9 
       (.I0(\stat_rd_data[30]_i_13_n_0 ),
        .I1(\stat_rd_data[30]_i_14_n_0 ),
        .O(\stat_rd_data_reg[30]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[31] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[31]),
        .Q(stat_rd_data[31]));
  MUXF8 \stat_rd_data_reg[31]_i_4 
       (.I0(\stat_rd_data_reg[31]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[31]_i_9_n_0 ),
        .O(\stat_rd_data_reg[31]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[31]_i_8 
       (.I0(\stat_rd_data[31]_i_11_n_0 ),
        .I1(\stat_rd_data[31]_i_12_n_0 ),
        .O(\stat_rd_data_reg[31]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[31]_i_9 
       (.I0(\stat_rd_data[31]_i_13_n_0 ),
        .I1(\stat_rd_data[31]_i_14_n_0 ),
        .O(\stat_rd_data_reg[31]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[32] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[32]),
        .Q(stat_rd_data[32]));
  MUXF8 \stat_rd_data_reg[32]_i_4 
       (.I0(\stat_rd_data_reg[32]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[32]_i_9_n_0 ),
        .O(\stat_rd_data_reg[32]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[32]_i_8 
       (.I0(\stat_rd_data[32]_i_11_n_0 ),
        .I1(\stat_rd_data[32]_i_12_n_0 ),
        .O(\stat_rd_data_reg[32]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[32]_i_9 
       (.I0(\stat_rd_data[32]_i_13_n_0 ),
        .I1(\stat_rd_data[32]_i_14_n_0 ),
        .O(\stat_rd_data_reg[32]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[33] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[33]),
        .Q(stat_rd_data[33]));
  MUXF8 \stat_rd_data_reg[33]_i_4 
       (.I0(\stat_rd_data_reg[33]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[33]_i_9_n_0 ),
        .O(\stat_rd_data_reg[33]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[33]_i_8 
       (.I0(\stat_rd_data[33]_i_11_n_0 ),
        .I1(\stat_rd_data[33]_i_12_n_0 ),
        .O(\stat_rd_data_reg[33]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[33]_i_9 
       (.I0(\stat_rd_data[33]_i_13_n_0 ),
        .I1(\stat_rd_data[33]_i_14_n_0 ),
        .O(\stat_rd_data_reg[33]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[34] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[34]),
        .Q(stat_rd_data[34]));
  MUXF8 \stat_rd_data_reg[34]_i_4 
       (.I0(\stat_rd_data_reg[34]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[34]_i_9_n_0 ),
        .O(\stat_rd_data_reg[34]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[34]_i_8 
       (.I0(\stat_rd_data[34]_i_11_n_0 ),
        .I1(\stat_rd_data[34]_i_12_n_0 ),
        .O(\stat_rd_data_reg[34]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[34]_i_9 
       (.I0(\stat_rd_data[34]_i_13_n_0 ),
        .I1(\stat_rd_data[34]_i_14_n_0 ),
        .O(\stat_rd_data_reg[34]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[35] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[35]),
        .Q(stat_rd_data[35]));
  MUXF8 \stat_rd_data_reg[35]_i_4 
       (.I0(\stat_rd_data_reg[35]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[35]_i_9_n_0 ),
        .O(\stat_rd_data_reg[35]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[35]_i_8 
       (.I0(\stat_rd_data[35]_i_11_n_0 ),
        .I1(\stat_rd_data[35]_i_12_n_0 ),
        .O(\stat_rd_data_reg[35]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[35]_i_9 
       (.I0(\stat_rd_data[35]_i_13_n_0 ),
        .I1(\stat_rd_data[35]_i_14_n_0 ),
        .O(\stat_rd_data_reg[35]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[36] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[36]),
        .Q(stat_rd_data[36]));
  MUXF8 \stat_rd_data_reg[36]_i_4 
       (.I0(\stat_rd_data_reg[36]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[36]_i_9_n_0 ),
        .O(\stat_rd_data_reg[36]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[36]_i_8 
       (.I0(\stat_rd_data[36]_i_11_n_0 ),
        .I1(\stat_rd_data[36]_i_12_n_0 ),
        .O(\stat_rd_data_reg[36]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[36]_i_9 
       (.I0(\stat_rd_data[36]_i_13_n_0 ),
        .I1(\stat_rd_data[36]_i_14_n_0 ),
        .O(\stat_rd_data_reg[36]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[37] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[37]),
        .Q(stat_rd_data[37]));
  MUXF8 \stat_rd_data_reg[37]_i_4 
       (.I0(\stat_rd_data_reg[37]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[37]_i_9_n_0 ),
        .O(\stat_rd_data_reg[37]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[37]_i_8 
       (.I0(\stat_rd_data[37]_i_11_n_0 ),
        .I1(\stat_rd_data[37]_i_12_n_0 ),
        .O(\stat_rd_data_reg[37]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[37]_i_9 
       (.I0(\stat_rd_data[37]_i_13_n_0 ),
        .I1(\stat_rd_data[37]_i_14_n_0 ),
        .O(\stat_rd_data_reg[37]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[38] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[38]),
        .Q(stat_rd_data[38]));
  MUXF8 \stat_rd_data_reg[38]_i_4 
       (.I0(\stat_rd_data_reg[38]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[38]_i_9_n_0 ),
        .O(\stat_rd_data_reg[38]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[38]_i_8 
       (.I0(\stat_rd_data[38]_i_11_n_0 ),
        .I1(\stat_rd_data[38]_i_12_n_0 ),
        .O(\stat_rd_data_reg[38]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[38]_i_9 
       (.I0(\stat_rd_data[38]_i_13_n_0 ),
        .I1(\stat_rd_data[38]_i_14_n_0 ),
        .O(\stat_rd_data_reg[38]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[39] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[39]),
        .Q(stat_rd_data[39]));
  MUXF8 \stat_rd_data_reg[39]_i_4 
       (.I0(\stat_rd_data_reg[39]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[39]_i_9_n_0 ),
        .O(\stat_rd_data_reg[39]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[39]_i_8 
       (.I0(\stat_rd_data[39]_i_11_n_0 ),
        .I1(\stat_rd_data[39]_i_12_n_0 ),
        .O(\stat_rd_data_reg[39]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[39]_i_9 
       (.I0(\stat_rd_data[39]_i_13_n_0 ),
        .I1(\stat_rd_data[39]_i_14_n_0 ),
        .O(\stat_rd_data_reg[39]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[3] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[3]),
        .Q(stat_rd_data[3]));
  MUXF8 \stat_rd_data_reg[3]_i_4 
       (.I0(\stat_rd_data_reg[3]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[3]_i_9_n_0 ),
        .O(\stat_rd_data_reg[3]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[3]_i_8 
       (.I0(\stat_rd_data[3]_i_11_n_0 ),
        .I1(\stat_rd_data[3]_i_12_n_0 ),
        .O(\stat_rd_data_reg[3]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[3]_i_9 
       (.I0(\stat_rd_data[3]_i_13_n_0 ),
        .I1(\stat_rd_data[3]_i_14_n_0 ),
        .O(\stat_rd_data_reg[3]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[40] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[40]),
        .Q(stat_rd_data[40]));
  MUXF8 \stat_rd_data_reg[40]_i_4 
       (.I0(\stat_rd_data_reg[40]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[40]_i_9_n_0 ),
        .O(\stat_rd_data_reg[40]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[40]_i_8 
       (.I0(\stat_rd_data[40]_i_11_n_0 ),
        .I1(\stat_rd_data[40]_i_12_n_0 ),
        .O(\stat_rd_data_reg[40]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[40]_i_9 
       (.I0(\stat_rd_data[40]_i_13_n_0 ),
        .I1(\stat_rd_data[40]_i_14_n_0 ),
        .O(\stat_rd_data_reg[40]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[41] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[41]),
        .Q(stat_rd_data[41]));
  MUXF8 \stat_rd_data_reg[41]_i_4 
       (.I0(\stat_rd_data_reg[41]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[41]_i_9_n_0 ),
        .O(\stat_rd_data_reg[41]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[41]_i_8 
       (.I0(\stat_rd_data[41]_i_11_n_0 ),
        .I1(\stat_rd_data[41]_i_12_n_0 ),
        .O(\stat_rd_data_reg[41]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[41]_i_9 
       (.I0(\stat_rd_data[41]_i_13_n_0 ),
        .I1(\stat_rd_data[41]_i_14_n_0 ),
        .O(\stat_rd_data_reg[41]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[42] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[42]),
        .Q(stat_rd_data[42]));
  MUXF8 \stat_rd_data_reg[42]_i_4 
       (.I0(\stat_rd_data_reg[42]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[42]_i_9_n_0 ),
        .O(\stat_rd_data_reg[42]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[42]_i_8 
       (.I0(\stat_rd_data[42]_i_11_n_0 ),
        .I1(\stat_rd_data[42]_i_12_n_0 ),
        .O(\stat_rd_data_reg[42]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[42]_i_9 
       (.I0(\stat_rd_data[42]_i_13_n_0 ),
        .I1(\stat_rd_data[42]_i_14_n_0 ),
        .O(\stat_rd_data_reg[42]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[43] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[43]),
        .Q(stat_rd_data[43]));
  MUXF8 \stat_rd_data_reg[43]_i_4 
       (.I0(\stat_rd_data_reg[43]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[43]_i_9_n_0 ),
        .O(\stat_rd_data_reg[43]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[43]_i_8 
       (.I0(\stat_rd_data[43]_i_11_n_0 ),
        .I1(\stat_rd_data[43]_i_12_n_0 ),
        .O(\stat_rd_data_reg[43]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[43]_i_9 
       (.I0(\stat_rd_data[43]_i_13_n_0 ),
        .I1(\stat_rd_data[43]_i_14_n_0 ),
        .O(\stat_rd_data_reg[43]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[44] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[44]),
        .Q(stat_rd_data[44]));
  MUXF8 \stat_rd_data_reg[44]_i_4 
       (.I0(\stat_rd_data_reg[44]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[44]_i_9_n_0 ),
        .O(\stat_rd_data_reg[44]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[44]_i_8 
       (.I0(\stat_rd_data[44]_i_11_n_0 ),
        .I1(\stat_rd_data[44]_i_12_n_0 ),
        .O(\stat_rd_data_reg[44]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[44]_i_9 
       (.I0(\stat_rd_data[44]_i_13_n_0 ),
        .I1(\stat_rd_data[44]_i_14_n_0 ),
        .O(\stat_rd_data_reg[44]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[45] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[45]),
        .Q(stat_rd_data[45]));
  MUXF8 \stat_rd_data_reg[45]_i_4 
       (.I0(\stat_rd_data_reg[45]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[45]_i_9_n_0 ),
        .O(\stat_rd_data_reg[45]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[45]_i_8 
       (.I0(\stat_rd_data[45]_i_11_n_0 ),
        .I1(\stat_rd_data[45]_i_12_n_0 ),
        .O(\stat_rd_data_reg[45]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[45]_i_9 
       (.I0(\stat_rd_data[45]_i_13_n_0 ),
        .I1(\stat_rd_data[45]_i_14_n_0 ),
        .O(\stat_rd_data_reg[45]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[46] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[46]),
        .Q(stat_rd_data[46]));
  MUXF8 \stat_rd_data_reg[46]_i_4 
       (.I0(\stat_rd_data_reg[46]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[46]_i_9_n_0 ),
        .O(\stat_rd_data_reg[46]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[46]_i_8 
       (.I0(\stat_rd_data[46]_i_11_n_0 ),
        .I1(\stat_rd_data[46]_i_12_n_0 ),
        .O(\stat_rd_data_reg[46]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[46]_i_9 
       (.I0(\stat_rd_data[46]_i_13_n_0 ),
        .I1(\stat_rd_data[46]_i_14_n_0 ),
        .O(\stat_rd_data_reg[46]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[47] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[47]),
        .Q(stat_rd_data[47]));
  MUXF8 \stat_rd_data_reg[47]_i_4 
       (.I0(\stat_rd_data_reg[47]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[47]_i_9_n_0 ),
        .O(\stat_rd_data_reg[47]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[47]_i_8 
       (.I0(\stat_rd_data[47]_i_11_n_0 ),
        .I1(\stat_rd_data[47]_i_12_n_0 ),
        .O(\stat_rd_data_reg[47]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[47]_i_9 
       (.I0(\stat_rd_data[47]_i_13_n_0 ),
        .I1(\stat_rd_data[47]_i_14_n_0 ),
        .O(\stat_rd_data_reg[47]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[48] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[48]),
        .Q(stat_rd_data[48]));
  MUXF8 \stat_rd_data_reg[48]_i_4 
       (.I0(\stat_rd_data_reg[48]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[48]_i_9_n_0 ),
        .O(\stat_rd_data_reg[48]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[48]_i_8 
       (.I0(\stat_rd_data[48]_i_11_n_0 ),
        .I1(\stat_rd_data[48]_i_12_n_0 ),
        .O(\stat_rd_data_reg[48]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[48]_i_9 
       (.I0(\stat_rd_data[48]_i_13_n_0 ),
        .I1(\stat_rd_data[48]_i_14_n_0 ),
        .O(\stat_rd_data_reg[48]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[49] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[49]),
        .Q(stat_rd_data[49]));
  MUXF8 \stat_rd_data_reg[49]_i_4 
       (.I0(\stat_rd_data_reg[49]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[49]_i_9_n_0 ),
        .O(\stat_rd_data_reg[49]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[49]_i_8 
       (.I0(\stat_rd_data[49]_i_11_n_0 ),
        .I1(\stat_rd_data[49]_i_12_n_0 ),
        .O(\stat_rd_data_reg[49]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[49]_i_9 
       (.I0(\stat_rd_data[49]_i_13_n_0 ),
        .I1(\stat_rd_data[49]_i_14_n_0 ),
        .O(\stat_rd_data_reg[49]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[4] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[4]),
        .Q(stat_rd_data[4]));
  MUXF8 \stat_rd_data_reg[4]_i_4 
       (.I0(\stat_rd_data_reg[4]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[4]_i_9_n_0 ),
        .O(\stat_rd_data_reg[4]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[4]_i_8 
       (.I0(\stat_rd_data[4]_i_11_n_0 ),
        .I1(\stat_rd_data[4]_i_12_n_0 ),
        .O(\stat_rd_data_reg[4]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[4]_i_9 
       (.I0(\stat_rd_data[4]_i_13_n_0 ),
        .I1(\stat_rd_data[4]_i_14_n_0 ),
        .O(\stat_rd_data_reg[4]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[50] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[50]),
        .Q(stat_rd_data[50]));
  MUXF8 \stat_rd_data_reg[50]_i_4 
       (.I0(\stat_rd_data_reg[50]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[50]_i_9_n_0 ),
        .O(\stat_rd_data_reg[50]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[50]_i_8 
       (.I0(\stat_rd_data[50]_i_11_n_0 ),
        .I1(\stat_rd_data[50]_i_12_n_0 ),
        .O(\stat_rd_data_reg[50]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[50]_i_9 
       (.I0(\stat_rd_data[50]_i_13_n_0 ),
        .I1(\stat_rd_data[50]_i_14_n_0 ),
        .O(\stat_rd_data_reg[50]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[51] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[51]),
        .Q(stat_rd_data[51]));
  MUXF8 \stat_rd_data_reg[51]_i_4 
       (.I0(\stat_rd_data_reg[51]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[51]_i_9_n_0 ),
        .O(\stat_rd_data_reg[51]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[51]_i_8 
       (.I0(\stat_rd_data[51]_i_11_n_0 ),
        .I1(\stat_rd_data[51]_i_12_n_0 ),
        .O(\stat_rd_data_reg[51]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[51]_i_9 
       (.I0(\stat_rd_data[51]_i_13_n_0 ),
        .I1(\stat_rd_data[51]_i_14_n_0 ),
        .O(\stat_rd_data_reg[51]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[52] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[52]),
        .Q(stat_rd_data[52]));
  MUXF8 \stat_rd_data_reg[52]_i_4 
       (.I0(\stat_rd_data_reg[52]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[52]_i_9_n_0 ),
        .O(\stat_rd_data_reg[52]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[52]_i_8 
       (.I0(\stat_rd_data[52]_i_11_n_0 ),
        .I1(\stat_rd_data[52]_i_12_n_0 ),
        .O(\stat_rd_data_reg[52]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[52]_i_9 
       (.I0(\stat_rd_data[52]_i_13_n_0 ),
        .I1(\stat_rd_data[52]_i_14_n_0 ),
        .O(\stat_rd_data_reg[52]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[53] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[53]),
        .Q(stat_rd_data[53]));
  MUXF8 \stat_rd_data_reg[53]_i_4 
       (.I0(\stat_rd_data_reg[53]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[53]_i_9_n_0 ),
        .O(\stat_rd_data_reg[53]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[53]_i_8 
       (.I0(\stat_rd_data[53]_i_11_n_0 ),
        .I1(\stat_rd_data[53]_i_12_n_0 ),
        .O(\stat_rd_data_reg[53]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[53]_i_9 
       (.I0(\stat_rd_data[53]_i_13_n_0 ),
        .I1(\stat_rd_data[53]_i_14_n_0 ),
        .O(\stat_rd_data_reg[53]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[54] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[54]),
        .Q(stat_rd_data[54]));
  MUXF8 \stat_rd_data_reg[54]_i_4 
       (.I0(\stat_rd_data_reg[54]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[54]_i_9_n_0 ),
        .O(\stat_rd_data_reg[54]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[54]_i_8 
       (.I0(\stat_rd_data[54]_i_11_n_0 ),
        .I1(\stat_rd_data[54]_i_12_n_0 ),
        .O(\stat_rd_data_reg[54]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[54]_i_9 
       (.I0(\stat_rd_data[54]_i_13_n_0 ),
        .I1(\stat_rd_data[54]_i_14_n_0 ),
        .O(\stat_rd_data_reg[54]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[55] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[55]),
        .Q(stat_rd_data[55]));
  MUXF8 \stat_rd_data_reg[55]_i_4 
       (.I0(\stat_rd_data_reg[55]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[55]_i_9_n_0 ),
        .O(\stat_rd_data_reg[55]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[55]_i_8 
       (.I0(\stat_rd_data[55]_i_11_n_0 ),
        .I1(\stat_rd_data[55]_i_12_n_0 ),
        .O(\stat_rd_data_reg[55]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[55]_i_9 
       (.I0(\stat_rd_data[55]_i_13_n_0 ),
        .I1(\stat_rd_data[55]_i_14_n_0 ),
        .O(\stat_rd_data_reg[55]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[56] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[56]),
        .Q(stat_rd_data[56]));
  MUXF8 \stat_rd_data_reg[56]_i_4 
       (.I0(\stat_rd_data_reg[56]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[56]_i_9_n_0 ),
        .O(\stat_rd_data_reg[56]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[56]_i_8 
       (.I0(\stat_rd_data[56]_i_11_n_0 ),
        .I1(\stat_rd_data[56]_i_12_n_0 ),
        .O(\stat_rd_data_reg[56]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[56]_i_9 
       (.I0(\stat_rd_data[56]_i_13_n_0 ),
        .I1(\stat_rd_data[56]_i_14_n_0 ),
        .O(\stat_rd_data_reg[56]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[57] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[57]),
        .Q(stat_rd_data[57]));
  MUXF8 \stat_rd_data_reg[57]_i_4 
       (.I0(\stat_rd_data_reg[57]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[57]_i_9_n_0 ),
        .O(\stat_rd_data_reg[57]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[57]_i_8 
       (.I0(\stat_rd_data[57]_i_11_n_0 ),
        .I1(\stat_rd_data[57]_i_12_n_0 ),
        .O(\stat_rd_data_reg[57]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[57]_i_9 
       (.I0(\stat_rd_data[57]_i_13_n_0 ),
        .I1(\stat_rd_data[57]_i_14_n_0 ),
        .O(\stat_rd_data_reg[57]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[58] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[58]),
        .Q(stat_rd_data[58]));
  MUXF8 \stat_rd_data_reg[58]_i_4 
       (.I0(\stat_rd_data_reg[58]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[58]_i_9_n_0 ),
        .O(\stat_rd_data_reg[58]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[58]_i_8 
       (.I0(\stat_rd_data[58]_i_11_n_0 ),
        .I1(\stat_rd_data[58]_i_12_n_0 ),
        .O(\stat_rd_data_reg[58]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[58]_i_9 
       (.I0(\stat_rd_data[58]_i_13_n_0 ),
        .I1(\stat_rd_data[58]_i_14_n_0 ),
        .O(\stat_rd_data_reg[58]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[59] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[59]),
        .Q(stat_rd_data[59]));
  MUXF8 \stat_rd_data_reg[59]_i_4 
       (.I0(\stat_rd_data_reg[59]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[59]_i_9_n_0 ),
        .O(\stat_rd_data_reg[59]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[59]_i_8 
       (.I0(\stat_rd_data[59]_i_11_n_0 ),
        .I1(\stat_rd_data[59]_i_12_n_0 ),
        .O(\stat_rd_data_reg[59]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[59]_i_9 
       (.I0(\stat_rd_data[59]_i_13_n_0 ),
        .I1(\stat_rd_data[59]_i_14_n_0 ),
        .O(\stat_rd_data_reg[59]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[5] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[5]),
        .Q(stat_rd_data[5]));
  MUXF8 \stat_rd_data_reg[5]_i_4 
       (.I0(\stat_rd_data_reg[5]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[5]_i_9_n_0 ),
        .O(\stat_rd_data_reg[5]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[5]_i_8 
       (.I0(\stat_rd_data[5]_i_11_n_0 ),
        .I1(\stat_rd_data[5]_i_12_n_0 ),
        .O(\stat_rd_data_reg[5]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[5]_i_9 
       (.I0(\stat_rd_data[5]_i_13_n_0 ),
        .I1(\stat_rd_data[5]_i_14_n_0 ),
        .O(\stat_rd_data_reg[5]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[60] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[60]),
        .Q(stat_rd_data[60]));
  MUXF8 \stat_rd_data_reg[60]_i_4 
       (.I0(\stat_rd_data_reg[60]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[60]_i_9_n_0 ),
        .O(\stat_rd_data_reg[60]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[60]_i_8 
       (.I0(\stat_rd_data[60]_i_11_n_0 ),
        .I1(\stat_rd_data[60]_i_12_n_0 ),
        .O(\stat_rd_data_reg[60]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[60]_i_9 
       (.I0(\stat_rd_data[60]_i_13_n_0 ),
        .I1(\stat_rd_data[60]_i_14_n_0 ),
        .O(\stat_rd_data_reg[60]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[61] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[61]),
        .Q(stat_rd_data[61]));
  MUXF8 \stat_rd_data_reg[61]_i_4 
       (.I0(\stat_rd_data_reg[61]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[61]_i_9_n_0 ),
        .O(\stat_rd_data_reg[61]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[61]_i_8 
       (.I0(\stat_rd_data[61]_i_11_n_0 ),
        .I1(\stat_rd_data[61]_i_12_n_0 ),
        .O(\stat_rd_data_reg[61]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[61]_i_9 
       (.I0(\stat_rd_data[61]_i_13_n_0 ),
        .I1(\stat_rd_data[61]_i_14_n_0 ),
        .O(\stat_rd_data_reg[61]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[62] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[62]),
        .Q(stat_rd_data[62]));
  MUXF8 \stat_rd_data_reg[62]_i_4 
       (.I0(\stat_rd_data_reg[62]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[62]_i_9_n_0 ),
        .O(\stat_rd_data_reg[62]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[62]_i_8 
       (.I0(\stat_rd_data[62]_i_11_n_0 ),
        .I1(\stat_rd_data[62]_i_12_n_0 ),
        .O(\stat_rd_data_reg[62]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[62]_i_9 
       (.I0(\stat_rd_data[62]_i_13_n_0 ),
        .I1(\stat_rd_data[62]_i_14_n_0 ),
        .O(\stat_rd_data_reg[62]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[63] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[63]),
        .Q(stat_rd_data[63]));
  MUXF7 \stat_rd_data_reg[63]_i_14 
       (.I0(\stat_rd_data[63]_i_17_n_0 ),
        .I1(\stat_rd_data[63]_i_18_n_0 ),
        .O(\stat_rd_data_reg[63]_i_14_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[63]_i_15 
       (.I0(\stat_rd_data[63]_i_19_n_0 ),
        .I1(\stat_rd_data[63]_i_20_n_0 ),
        .O(\stat_rd_data_reg[63]_i_15_n_0 ),
        .S(out[2]));
  MUXF8 \stat_rd_data_reg[63]_i_8 
       (.I0(\stat_rd_data_reg[63]_i_14_n_0 ),
        .I1(\stat_rd_data_reg[63]_i_15_n_0 ),
        .O(\stat_rd_data_reg[63]_i_8_n_0 ),
        .S(out[3]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[6] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[6]),
        .Q(stat_rd_data[6]));
  MUXF8 \stat_rd_data_reg[6]_i_4 
       (.I0(\stat_rd_data_reg[6]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[6]_i_9_n_0 ),
        .O(\stat_rd_data_reg[6]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[6]_i_8 
       (.I0(\stat_rd_data[6]_i_11_n_0 ),
        .I1(\stat_rd_data[6]_i_12_n_0 ),
        .O(\stat_rd_data_reg[6]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[6]_i_9 
       (.I0(\stat_rd_data[6]_i_13_n_0 ),
        .I1(\stat_rd_data[6]_i_14_n_0 ),
        .O(\stat_rd_data_reg[6]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[7] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[7]),
        .Q(stat_rd_data[7]));
  MUXF8 \stat_rd_data_reg[7]_i_4 
       (.I0(\stat_rd_data_reg[7]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[7]_i_9_n_0 ),
        .O(\stat_rd_data_reg[7]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[7]_i_8 
       (.I0(\stat_rd_data[7]_i_11_n_0 ),
        .I1(\stat_rd_data[7]_i_12_n_0 ),
        .O(\stat_rd_data_reg[7]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[7]_i_9 
       (.I0(\stat_rd_data[7]_i_13_n_0 ),
        .I1(\stat_rd_data[7]_i_14_n_0 ),
        .O(\stat_rd_data_reg[7]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[8] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[8]),
        .Q(stat_rd_data[8]));
  MUXF8 \stat_rd_data_reg[8]_i_4 
       (.I0(\stat_rd_data_reg[8]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[8]_i_9_n_0 ),
        .O(\stat_rd_data_reg[8]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[8]_i_8 
       (.I0(\stat_rd_data[8]_i_11_n_0 ),
        .I1(\stat_rd_data[8]_i_12_n_0 ),
        .O(\stat_rd_data_reg[8]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[8]_i_9 
       (.I0(\stat_rd_data[8]_i_13_n_0 ),
        .I1(\stat_rd_data[8]_i_14_n_0 ),
        .O(\stat_rd_data_reg[8]_i_9_n_0 ),
        .S(out[2]));
  FDCE #(
    .INIT(1'b0)) 
    \stat_rd_data_reg[9] 
       (.C(clk_i),
        .CE(\stat_rd_data[63]_i_1_n_0 ),
        .CLR(rst_i),
        .D(p_0_in[9]),
        .Q(stat_rd_data[9]));
  MUXF8 \stat_rd_data_reg[9]_i_4 
       (.I0(\stat_rd_data_reg[9]_i_8_n_0 ),
        .I1(\stat_rd_data_reg[9]_i_9_n_0 ),
        .O(\stat_rd_data_reg[9]_i_4_n_0 ),
        .S(out[3]));
  MUXF7 \stat_rd_data_reg[9]_i_8 
       (.I0(\stat_rd_data[9]_i_11_n_0 ),
        .I1(\stat_rd_data[9]_i_12_n_0 ),
        .O(\stat_rd_data_reg[9]_i_8_n_0 ),
        .S(out[2]));
  MUXF7 \stat_rd_data_reg[9]_i_9 
       (.I0(\stat_rd_data[9]_i_13_n_0 ),
        .I1(\stat_rd_data[9]_i_14_n_0 ),
        .O(\stat_rd_data_reg[9]_i_9_n_0 ),
        .S(out[2]));
  LUT6 #(
    .INIT(64'hCC0CC00077477444)) 
    \state[0]_i_1 
       (.I0(state1__0),
        .I1(\state_reg_n_0_[0] ),
        .I2(\stat_rd_data_reg[63]_1 ),
        .I3(\stat_rd_data_reg[63]_0 ),
        .I4(out[9]),
        .I5(\state_reg_n_0_[1] ),
        .O(state[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \state[0]_i_2 
       (.I0(mdio_in_valid_d1),
        .I1(mdio_in_valid),
        .O(state1__0));
  LUT6 #(
    .INIT(64'h1010B5B51010B510)) 
    \state[1]_i_1 
       (.I0(\state_reg_n_0_[0] ),
        .I1(read_done_reg_n_0),
        .I2(\state_reg_n_0_[1] ),
        .I3(out[9]),
        .I4(\stat_rd_data_reg[63]_1 ),
        .I5(\stat_rd_data_reg[63]_0 ),
        .O(state[1]));
  FDCE #(
    .INIT(1'b0)) 
    \state_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(state[0]),
        .Q(\state_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \state_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(state[1]),
        .Q(\state_reg_n_0_[1] ));
  LUT1 #(
    .INIT(2'h1)) 
    \tagged_frame_good[0]_i_2 
       (.I0(tagged_frame_good_reg[0]),
        .O(\tagged_frame_good[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[0]_i_1_n_0 ,\tagged_frame_good_reg[0]_i_1_n_1 ,\tagged_frame_good_reg[0]_i_1_n_2 ,\tagged_frame_good_reg[0]_i_1_n_3 ,\tagged_frame_good_reg[0]_i_1_n_4 ,\tagged_frame_good_reg[0]_i_1_n_5 ,\tagged_frame_good_reg[0]_i_1_n_6 ,\tagged_frame_good_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\tagged_frame_good_reg[0]_i_1_n_8 ,\tagged_frame_good_reg[0]_i_1_n_9 ,\tagged_frame_good_reg[0]_i_1_n_10 ,\tagged_frame_good_reg[0]_i_1_n_11 ,\tagged_frame_good_reg[0]_i_1_n_12 ,\tagged_frame_good_reg[0]_i_1_n_13 ,\tagged_frame_good_reg[0]_i_1_n_14 ,\tagged_frame_good_reg[0]_i_1_n_15 }),
        .S({tagged_frame_good_reg[7:1],\tagged_frame_good[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[16]_i_1 
       (.CI(\tagged_frame_good_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[16]_i_1_n_0 ,\tagged_frame_good_reg[16]_i_1_n_1 ,\tagged_frame_good_reg[16]_i_1_n_2 ,\tagged_frame_good_reg[16]_i_1_n_3 ,\tagged_frame_good_reg[16]_i_1_n_4 ,\tagged_frame_good_reg[16]_i_1_n_5 ,\tagged_frame_good_reg[16]_i_1_n_6 ,\tagged_frame_good_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[16]_i_1_n_8 ,\tagged_frame_good_reg[16]_i_1_n_9 ,\tagged_frame_good_reg[16]_i_1_n_10 ,\tagged_frame_good_reg[16]_i_1_n_11 ,\tagged_frame_good_reg[16]_i_1_n_12 ,\tagged_frame_good_reg[16]_i_1_n_13 ,\tagged_frame_good_reg[16]_i_1_n_14 ,\tagged_frame_good_reg[16]_i_1_n_15 }),
        .S(tagged_frame_good_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[16]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[24]_i_1 
       (.CI(\tagged_frame_good_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[24]_i_1_n_0 ,\tagged_frame_good_reg[24]_i_1_n_1 ,\tagged_frame_good_reg[24]_i_1_n_2 ,\tagged_frame_good_reg[24]_i_1_n_3 ,\tagged_frame_good_reg[24]_i_1_n_4 ,\tagged_frame_good_reg[24]_i_1_n_5 ,\tagged_frame_good_reg[24]_i_1_n_6 ,\tagged_frame_good_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[24]_i_1_n_8 ,\tagged_frame_good_reg[24]_i_1_n_9 ,\tagged_frame_good_reg[24]_i_1_n_10 ,\tagged_frame_good_reg[24]_i_1_n_11 ,\tagged_frame_good_reg[24]_i_1_n_12 ,\tagged_frame_good_reg[24]_i_1_n_13 ,\tagged_frame_good_reg[24]_i_1_n_14 ,\tagged_frame_good_reg[24]_i_1_n_15 }),
        .S(tagged_frame_good_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[24]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[32]_i_1 
       (.CI(\tagged_frame_good_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[32]_i_1_n_0 ,\tagged_frame_good_reg[32]_i_1_n_1 ,\tagged_frame_good_reg[32]_i_1_n_2 ,\tagged_frame_good_reg[32]_i_1_n_3 ,\tagged_frame_good_reg[32]_i_1_n_4 ,\tagged_frame_good_reg[32]_i_1_n_5 ,\tagged_frame_good_reg[32]_i_1_n_6 ,\tagged_frame_good_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[32]_i_1_n_8 ,\tagged_frame_good_reg[32]_i_1_n_9 ,\tagged_frame_good_reg[32]_i_1_n_10 ,\tagged_frame_good_reg[32]_i_1_n_11 ,\tagged_frame_good_reg[32]_i_1_n_12 ,\tagged_frame_good_reg[32]_i_1_n_13 ,\tagged_frame_good_reg[32]_i_1_n_14 ,\tagged_frame_good_reg[32]_i_1_n_15 }),
        .S(tagged_frame_good_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[32]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[40]_i_1 
       (.CI(\tagged_frame_good_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[40]_i_1_n_0 ,\tagged_frame_good_reg[40]_i_1_n_1 ,\tagged_frame_good_reg[40]_i_1_n_2 ,\tagged_frame_good_reg[40]_i_1_n_3 ,\tagged_frame_good_reg[40]_i_1_n_4 ,\tagged_frame_good_reg[40]_i_1_n_5 ,\tagged_frame_good_reg[40]_i_1_n_6 ,\tagged_frame_good_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[40]_i_1_n_8 ,\tagged_frame_good_reg[40]_i_1_n_9 ,\tagged_frame_good_reg[40]_i_1_n_10 ,\tagged_frame_good_reg[40]_i_1_n_11 ,\tagged_frame_good_reg[40]_i_1_n_12 ,\tagged_frame_good_reg[40]_i_1_n_13 ,\tagged_frame_good_reg[40]_i_1_n_14 ,\tagged_frame_good_reg[40]_i_1_n_15 }),
        .S(tagged_frame_good_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[40]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[48]_i_1 
       (.CI(\tagged_frame_good_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[48]_i_1_n_0 ,\tagged_frame_good_reg[48]_i_1_n_1 ,\tagged_frame_good_reg[48]_i_1_n_2 ,\tagged_frame_good_reg[48]_i_1_n_3 ,\tagged_frame_good_reg[48]_i_1_n_4 ,\tagged_frame_good_reg[48]_i_1_n_5 ,\tagged_frame_good_reg[48]_i_1_n_6 ,\tagged_frame_good_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[48]_i_1_n_8 ,\tagged_frame_good_reg[48]_i_1_n_9 ,\tagged_frame_good_reg[48]_i_1_n_10 ,\tagged_frame_good_reg[48]_i_1_n_11 ,\tagged_frame_good_reg[48]_i_1_n_12 ,\tagged_frame_good_reg[48]_i_1_n_13 ,\tagged_frame_good_reg[48]_i_1_n_14 ,\tagged_frame_good_reg[48]_i_1_n_15 }),
        .S(tagged_frame_good_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[48]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[56]_i_1 
       (.CI(\tagged_frame_good_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_tagged_frame_good_reg[56]_i_1_CO_UNCONNECTED [7],\tagged_frame_good_reg[56]_i_1_n_1 ,\tagged_frame_good_reg[56]_i_1_n_2 ,\tagged_frame_good_reg[56]_i_1_n_3 ,\tagged_frame_good_reg[56]_i_1_n_4 ,\tagged_frame_good_reg[56]_i_1_n_5 ,\tagged_frame_good_reg[56]_i_1_n_6 ,\tagged_frame_good_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[56]_i_1_n_8 ,\tagged_frame_good_reg[56]_i_1_n_9 ,\tagged_frame_good_reg[56]_i_1_n_10 ,\tagged_frame_good_reg[56]_i_1_n_11 ,\tagged_frame_good_reg[56]_i_1_n_12 ,\tagged_frame_good_reg[56]_i_1_n_13 ,\tagged_frame_good_reg[56]_i_1_n_14 ,\tagged_frame_good_reg[56]_i_1_n_15 }),
        .S(tagged_frame_good_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_13 ),
        .Q(tagged_frame_good_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_12 ),
        .Q(tagged_frame_good_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_11 ),
        .Q(tagged_frame_good_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_10 ),
        .Q(tagged_frame_good_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[56]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_9 ),
        .Q(tagged_frame_good_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[0]_i_1_n_8 ),
        .Q(tagged_frame_good_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_15 ),
        .Q(tagged_frame_good_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_good_reg[8]_i_1 
       (.CI(\tagged_frame_good_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_good_reg[8]_i_1_n_0 ,\tagged_frame_good_reg[8]_i_1_n_1 ,\tagged_frame_good_reg[8]_i_1_n_2 ,\tagged_frame_good_reg[8]_i_1_n_3 ,\tagged_frame_good_reg[8]_i_1_n_4 ,\tagged_frame_good_reg[8]_i_1_n_5 ,\tagged_frame_good_reg[8]_i_1_n_6 ,\tagged_frame_good_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_good_reg[8]_i_1_n_8 ,\tagged_frame_good_reg[8]_i_1_n_9 ,\tagged_frame_good_reg[8]_i_1_n_10 ,\tagged_frame_good_reg[8]_i_1_n_11 ,\tagged_frame_good_reg[8]_i_1_n_12 ,\tagged_frame_good_reg[8]_i_1_n_13 ,\tagged_frame_good_reg[8]_i_1_n_14 ,\tagged_frame_good_reg[8]_i_1_n_15 }),
        .S(tagged_frame_good_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_good_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_good_reg[8]_i_1_n_14 ),
        .Q(tagged_frame_good_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \tagged_frame_transed[0]_i_2 
       (.I0(tagged_frame_transed_reg[0]),
        .O(\tagged_frame_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[0]_i_1_n_0 ,\tagged_frame_transed_reg[0]_i_1_n_1 ,\tagged_frame_transed_reg[0]_i_1_n_2 ,\tagged_frame_transed_reg[0]_i_1_n_3 ,\tagged_frame_transed_reg[0]_i_1_n_4 ,\tagged_frame_transed_reg[0]_i_1_n_5 ,\tagged_frame_transed_reg[0]_i_1_n_6 ,\tagged_frame_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\tagged_frame_transed_reg[0]_i_1_n_8 ,\tagged_frame_transed_reg[0]_i_1_n_9 ,\tagged_frame_transed_reg[0]_i_1_n_10 ,\tagged_frame_transed_reg[0]_i_1_n_11 ,\tagged_frame_transed_reg[0]_i_1_n_12 ,\tagged_frame_transed_reg[0]_i_1_n_13 ,\tagged_frame_transed_reg[0]_i_1_n_14 ,\tagged_frame_transed_reg[0]_i_1_n_15 }),
        .S({tagged_frame_transed_reg[7:1],\tagged_frame_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[16]_i_1 
       (.CI(\tagged_frame_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[16]_i_1_n_0 ,\tagged_frame_transed_reg[16]_i_1_n_1 ,\tagged_frame_transed_reg[16]_i_1_n_2 ,\tagged_frame_transed_reg[16]_i_1_n_3 ,\tagged_frame_transed_reg[16]_i_1_n_4 ,\tagged_frame_transed_reg[16]_i_1_n_5 ,\tagged_frame_transed_reg[16]_i_1_n_6 ,\tagged_frame_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[16]_i_1_n_8 ,\tagged_frame_transed_reg[16]_i_1_n_9 ,\tagged_frame_transed_reg[16]_i_1_n_10 ,\tagged_frame_transed_reg[16]_i_1_n_11 ,\tagged_frame_transed_reg[16]_i_1_n_12 ,\tagged_frame_transed_reg[16]_i_1_n_13 ,\tagged_frame_transed_reg[16]_i_1_n_14 ,\tagged_frame_transed_reg[16]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[16]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[24]_i_1 
       (.CI(\tagged_frame_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[24]_i_1_n_0 ,\tagged_frame_transed_reg[24]_i_1_n_1 ,\tagged_frame_transed_reg[24]_i_1_n_2 ,\tagged_frame_transed_reg[24]_i_1_n_3 ,\tagged_frame_transed_reg[24]_i_1_n_4 ,\tagged_frame_transed_reg[24]_i_1_n_5 ,\tagged_frame_transed_reg[24]_i_1_n_6 ,\tagged_frame_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[24]_i_1_n_8 ,\tagged_frame_transed_reg[24]_i_1_n_9 ,\tagged_frame_transed_reg[24]_i_1_n_10 ,\tagged_frame_transed_reg[24]_i_1_n_11 ,\tagged_frame_transed_reg[24]_i_1_n_12 ,\tagged_frame_transed_reg[24]_i_1_n_13 ,\tagged_frame_transed_reg[24]_i_1_n_14 ,\tagged_frame_transed_reg[24]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[24]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[32]_i_1 
       (.CI(\tagged_frame_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[32]_i_1_n_0 ,\tagged_frame_transed_reg[32]_i_1_n_1 ,\tagged_frame_transed_reg[32]_i_1_n_2 ,\tagged_frame_transed_reg[32]_i_1_n_3 ,\tagged_frame_transed_reg[32]_i_1_n_4 ,\tagged_frame_transed_reg[32]_i_1_n_5 ,\tagged_frame_transed_reg[32]_i_1_n_6 ,\tagged_frame_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[32]_i_1_n_8 ,\tagged_frame_transed_reg[32]_i_1_n_9 ,\tagged_frame_transed_reg[32]_i_1_n_10 ,\tagged_frame_transed_reg[32]_i_1_n_11 ,\tagged_frame_transed_reg[32]_i_1_n_12 ,\tagged_frame_transed_reg[32]_i_1_n_13 ,\tagged_frame_transed_reg[32]_i_1_n_14 ,\tagged_frame_transed_reg[32]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[32]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[40]_i_1 
       (.CI(\tagged_frame_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[40]_i_1_n_0 ,\tagged_frame_transed_reg[40]_i_1_n_1 ,\tagged_frame_transed_reg[40]_i_1_n_2 ,\tagged_frame_transed_reg[40]_i_1_n_3 ,\tagged_frame_transed_reg[40]_i_1_n_4 ,\tagged_frame_transed_reg[40]_i_1_n_5 ,\tagged_frame_transed_reg[40]_i_1_n_6 ,\tagged_frame_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[40]_i_1_n_8 ,\tagged_frame_transed_reg[40]_i_1_n_9 ,\tagged_frame_transed_reg[40]_i_1_n_10 ,\tagged_frame_transed_reg[40]_i_1_n_11 ,\tagged_frame_transed_reg[40]_i_1_n_12 ,\tagged_frame_transed_reg[40]_i_1_n_13 ,\tagged_frame_transed_reg[40]_i_1_n_14 ,\tagged_frame_transed_reg[40]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[40]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[48]_i_1 
       (.CI(\tagged_frame_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[48]_i_1_n_0 ,\tagged_frame_transed_reg[48]_i_1_n_1 ,\tagged_frame_transed_reg[48]_i_1_n_2 ,\tagged_frame_transed_reg[48]_i_1_n_3 ,\tagged_frame_transed_reg[48]_i_1_n_4 ,\tagged_frame_transed_reg[48]_i_1_n_5 ,\tagged_frame_transed_reg[48]_i_1_n_6 ,\tagged_frame_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[48]_i_1_n_8 ,\tagged_frame_transed_reg[48]_i_1_n_9 ,\tagged_frame_transed_reg[48]_i_1_n_10 ,\tagged_frame_transed_reg[48]_i_1_n_11 ,\tagged_frame_transed_reg[48]_i_1_n_12 ,\tagged_frame_transed_reg[48]_i_1_n_13 ,\tagged_frame_transed_reg[48]_i_1_n_14 ,\tagged_frame_transed_reg[48]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[48]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[56]_i_1 
       (.CI(\tagged_frame_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_tagged_frame_transed_reg[56]_i_1_CO_UNCONNECTED [7],\tagged_frame_transed_reg[56]_i_1_n_1 ,\tagged_frame_transed_reg[56]_i_1_n_2 ,\tagged_frame_transed_reg[56]_i_1_n_3 ,\tagged_frame_transed_reg[56]_i_1_n_4 ,\tagged_frame_transed_reg[56]_i_1_n_5 ,\tagged_frame_transed_reg[56]_i_1_n_6 ,\tagged_frame_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[56]_i_1_n_8 ,\tagged_frame_transed_reg[56]_i_1_n_9 ,\tagged_frame_transed_reg[56]_i_1_n_10 ,\tagged_frame_transed_reg[56]_i_1_n_11 ,\tagged_frame_transed_reg[56]_i_1_n_12 ,\tagged_frame_transed_reg[56]_i_1_n_13 ,\tagged_frame_transed_reg[56]_i_1_n_14 ,\tagged_frame_transed_reg[56]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_13 ),
        .Q(tagged_frame_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_12 ),
        .Q(tagged_frame_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_11 ),
        .Q(tagged_frame_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_10 ),
        .Q(tagged_frame_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[56]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_9 ),
        .Q(tagged_frame_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[0]_i_1_n_8 ),
        .Q(tagged_frame_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_15 ),
        .Q(tagged_frame_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \tagged_frame_transed_reg[8]_i_1 
       (.CI(\tagged_frame_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\tagged_frame_transed_reg[8]_i_1_n_0 ,\tagged_frame_transed_reg[8]_i_1_n_1 ,\tagged_frame_transed_reg[8]_i_1_n_2 ,\tagged_frame_transed_reg[8]_i_1_n_3 ,\tagged_frame_transed_reg[8]_i_1_n_4 ,\tagged_frame_transed_reg[8]_i_1_n_5 ,\tagged_frame_transed_reg[8]_i_1_n_6 ,\tagged_frame_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\tagged_frame_transed_reg[8]_i_1_n_8 ,\tagged_frame_transed_reg[8]_i_1_n_9 ,\tagged_frame_transed_reg[8]_i_1_n_10 ,\tagged_frame_transed_reg[8]_i_1_n_11 ,\tagged_frame_transed_reg[8]_i_1_n_12 ,\tagged_frame_transed_reg[8]_i_1_n_13 ,\tagged_frame_transed_reg[8]_i_1_n_14 ,\tagged_frame_transed_reg[8]_i_1_n_15 }),
        .S(tagged_frame_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \tagged_frame_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[12]),
        .CLR(rst_i),
        .D(\tagged_frame_transed_reg[8]_i_1_n_14 ),
        .Q(tagged_frame_transed_reg[9]));
  LUT6 #(
    .INIT(64'h0000000015555555)) 
    \tmp_cnt[0]_i_1 
       (.I0(tmp_cnt[0]),
        .I1(tmp_cnt[2]),
        .I2(tmp_cnt[1]),
        .I3(tmp_cnt[3]),
        .I4(tmp_cnt[4]),
        .I5(state15_out),
        .O(\tmp_cnt[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \tmp_cnt[1]_i_1 
       (.I0(tmp_cnt[0]),
        .I1(tmp_cnt[1]),
        .I2(state15_out),
        .O(\tmp_cnt[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT4 #(
    .INIT(16'h0078)) 
    \tmp_cnt[2]_i_1 
       (.I0(tmp_cnt[0]),
        .I1(tmp_cnt[1]),
        .I2(tmp_cnt[2]),
        .I3(state15_out),
        .O(\tmp_cnt[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT5 #(
    .INIT(32'h000078F0)) 
    \tmp_cnt[3]_i_1 
       (.I0(tmp_cnt[0]),
        .I1(tmp_cnt[1]),
        .I2(tmp_cnt[3]),
        .I3(tmp_cnt[2]),
        .I4(state15_out),
        .O(\tmp_cnt[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000078F0F0F0)) 
    \tmp_cnt[4]_i_1 
       (.I0(tmp_cnt[0]),
        .I1(tmp_cnt[1]),
        .I2(tmp_cnt[4]),
        .I3(tmp_cnt[3]),
        .I4(tmp_cnt[2]),
        .I5(state15_out),
        .O(\tmp_cnt[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \tmp_cnt[4]_i_2 
       (.I0(\stat_rd_data_reg[63]_0 ),
        .I1(\stat_rd_data_reg[63]_1 ),
        .O(state15_out));
  FDCE #(
    .INIT(1'b0)) 
    \tmp_cnt_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\tmp_cnt[0]_i_1_n_0 ),
        .Q(tmp_cnt[0]));
  FDCE #(
    .INIT(1'b0)) 
    \tmp_cnt_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\tmp_cnt[1]_i_1_n_0 ),
        .Q(tmp_cnt[1]));
  FDCE #(
    .INIT(1'b0)) 
    \tmp_cnt_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\tmp_cnt[2]_i_1_n_0 ),
        .Q(tmp_cnt[2]));
  FDCE #(
    .INIT(1'b0)) 
    \tmp_cnt_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\tmp_cnt[3]_i_1_n_0 ),
        .Q(tmp_cnt[3]));
  FDCE #(
    .INIT(1'b0)) 
    \tmp_cnt_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\tmp_cnt[4]_i_1_n_0 ),
        .Q(tmp_cnt[4]));
  LUT1 #(
    .INIT(2'h1)) 
    \total_bytes_recved[0]_i_2 
       (.I0(total_bytes_recved_reg[0]),
        .O(\total_bytes_recved[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[0]_i_1_n_0 ,\total_bytes_recved_reg[0]_i_1_n_1 ,\total_bytes_recved_reg[0]_i_1_n_2 ,\total_bytes_recved_reg[0]_i_1_n_3 ,\total_bytes_recved_reg[0]_i_1_n_4 ,\total_bytes_recved_reg[0]_i_1_n_5 ,\total_bytes_recved_reg[0]_i_1_n_6 ,\total_bytes_recved_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\total_bytes_recved_reg[0]_i_1_n_8 ,\total_bytes_recved_reg[0]_i_1_n_9 ,\total_bytes_recved_reg[0]_i_1_n_10 ,\total_bytes_recved_reg[0]_i_1_n_11 ,\total_bytes_recved_reg[0]_i_1_n_12 ,\total_bytes_recved_reg[0]_i_1_n_13 ,\total_bytes_recved_reg[0]_i_1_n_14 ,\total_bytes_recved_reg[0]_i_1_n_15 }),
        .S({total_bytes_recved_reg[7:1],\total_bytes_recved[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[16]_i_1 
       (.CI(\total_bytes_recved_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[16]_i_1_n_0 ,\total_bytes_recved_reg[16]_i_1_n_1 ,\total_bytes_recved_reg[16]_i_1_n_2 ,\total_bytes_recved_reg[16]_i_1_n_3 ,\total_bytes_recved_reg[16]_i_1_n_4 ,\total_bytes_recved_reg[16]_i_1_n_5 ,\total_bytes_recved_reg[16]_i_1_n_6 ,\total_bytes_recved_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[16]_i_1_n_8 ,\total_bytes_recved_reg[16]_i_1_n_9 ,\total_bytes_recved_reg[16]_i_1_n_10 ,\total_bytes_recved_reg[16]_i_1_n_11 ,\total_bytes_recved_reg[16]_i_1_n_12 ,\total_bytes_recved_reg[16]_i_1_n_13 ,\total_bytes_recved_reg[16]_i_1_n_14 ,\total_bytes_recved_reg[16]_i_1_n_15 }),
        .S(total_bytes_recved_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[16]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[24]_i_1 
       (.CI(\total_bytes_recved_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[24]_i_1_n_0 ,\total_bytes_recved_reg[24]_i_1_n_1 ,\total_bytes_recved_reg[24]_i_1_n_2 ,\total_bytes_recved_reg[24]_i_1_n_3 ,\total_bytes_recved_reg[24]_i_1_n_4 ,\total_bytes_recved_reg[24]_i_1_n_5 ,\total_bytes_recved_reg[24]_i_1_n_6 ,\total_bytes_recved_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[24]_i_1_n_8 ,\total_bytes_recved_reg[24]_i_1_n_9 ,\total_bytes_recved_reg[24]_i_1_n_10 ,\total_bytes_recved_reg[24]_i_1_n_11 ,\total_bytes_recved_reg[24]_i_1_n_12 ,\total_bytes_recved_reg[24]_i_1_n_13 ,\total_bytes_recved_reg[24]_i_1_n_14 ,\total_bytes_recved_reg[24]_i_1_n_15 }),
        .S(total_bytes_recved_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[24]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[32]_i_1 
       (.CI(\total_bytes_recved_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[32]_i_1_n_0 ,\total_bytes_recved_reg[32]_i_1_n_1 ,\total_bytes_recved_reg[32]_i_1_n_2 ,\total_bytes_recved_reg[32]_i_1_n_3 ,\total_bytes_recved_reg[32]_i_1_n_4 ,\total_bytes_recved_reg[32]_i_1_n_5 ,\total_bytes_recved_reg[32]_i_1_n_6 ,\total_bytes_recved_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[32]_i_1_n_8 ,\total_bytes_recved_reg[32]_i_1_n_9 ,\total_bytes_recved_reg[32]_i_1_n_10 ,\total_bytes_recved_reg[32]_i_1_n_11 ,\total_bytes_recved_reg[32]_i_1_n_12 ,\total_bytes_recved_reg[32]_i_1_n_13 ,\total_bytes_recved_reg[32]_i_1_n_14 ,\total_bytes_recved_reg[32]_i_1_n_15 }),
        .S(total_bytes_recved_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[32]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[40]_i_1 
       (.CI(\total_bytes_recved_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[40]_i_1_n_0 ,\total_bytes_recved_reg[40]_i_1_n_1 ,\total_bytes_recved_reg[40]_i_1_n_2 ,\total_bytes_recved_reg[40]_i_1_n_3 ,\total_bytes_recved_reg[40]_i_1_n_4 ,\total_bytes_recved_reg[40]_i_1_n_5 ,\total_bytes_recved_reg[40]_i_1_n_6 ,\total_bytes_recved_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[40]_i_1_n_8 ,\total_bytes_recved_reg[40]_i_1_n_9 ,\total_bytes_recved_reg[40]_i_1_n_10 ,\total_bytes_recved_reg[40]_i_1_n_11 ,\total_bytes_recved_reg[40]_i_1_n_12 ,\total_bytes_recved_reg[40]_i_1_n_13 ,\total_bytes_recved_reg[40]_i_1_n_14 ,\total_bytes_recved_reg[40]_i_1_n_15 }),
        .S(total_bytes_recved_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[40]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[48]_i_1 
       (.CI(\total_bytes_recved_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[48]_i_1_n_0 ,\total_bytes_recved_reg[48]_i_1_n_1 ,\total_bytes_recved_reg[48]_i_1_n_2 ,\total_bytes_recved_reg[48]_i_1_n_3 ,\total_bytes_recved_reg[48]_i_1_n_4 ,\total_bytes_recved_reg[48]_i_1_n_5 ,\total_bytes_recved_reg[48]_i_1_n_6 ,\total_bytes_recved_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[48]_i_1_n_8 ,\total_bytes_recved_reg[48]_i_1_n_9 ,\total_bytes_recved_reg[48]_i_1_n_10 ,\total_bytes_recved_reg[48]_i_1_n_11 ,\total_bytes_recved_reg[48]_i_1_n_12 ,\total_bytes_recved_reg[48]_i_1_n_13 ,\total_bytes_recved_reg[48]_i_1_n_14 ,\total_bytes_recved_reg[48]_i_1_n_15 }),
        .S(total_bytes_recved_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[48]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[56]_i_1 
       (.CI(\total_bytes_recved_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_total_bytes_recved_reg[56]_i_1_CO_UNCONNECTED [7],\total_bytes_recved_reg[56]_i_1_n_1 ,\total_bytes_recved_reg[56]_i_1_n_2 ,\total_bytes_recved_reg[56]_i_1_n_3 ,\total_bytes_recved_reg[56]_i_1_n_4 ,\total_bytes_recved_reg[56]_i_1_n_5 ,\total_bytes_recved_reg[56]_i_1_n_6 ,\total_bytes_recved_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[56]_i_1_n_8 ,\total_bytes_recved_reg[56]_i_1_n_9 ,\total_bytes_recved_reg[56]_i_1_n_10 ,\total_bytes_recved_reg[56]_i_1_n_11 ,\total_bytes_recved_reg[56]_i_1_n_12 ,\total_bytes_recved_reg[56]_i_1_n_13 ,\total_bytes_recved_reg[56]_i_1_n_14 ,\total_bytes_recved_reg[56]_i_1_n_15 }),
        .S(total_bytes_recved_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_13 ),
        .Q(total_bytes_recved_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_12 ),
        .Q(total_bytes_recved_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_11 ),
        .Q(total_bytes_recved_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_10 ),
        .Q(total_bytes_recved_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[56]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_9 ),
        .Q(total_bytes_recved_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[0]_i_1_n_8 ),
        .Q(total_bytes_recved_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_15 ),
        .Q(total_bytes_recved_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_recved_reg[8]_i_1 
       (.CI(\total_bytes_recved_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_recved_reg[8]_i_1_n_0 ,\total_bytes_recved_reg[8]_i_1_n_1 ,\total_bytes_recved_reg[8]_i_1_n_2 ,\total_bytes_recved_reg[8]_i_1_n_3 ,\total_bytes_recved_reg[8]_i_1_n_4 ,\total_bytes_recved_reg[8]_i_1_n_5 ,\total_bytes_recved_reg[8]_i_1_n_6 ,\total_bytes_recved_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_recved_reg[8]_i_1_n_8 ,\total_bytes_recved_reg[8]_i_1_n_9 ,\total_bytes_recved_reg[8]_i_1_n_10 ,\total_bytes_recved_reg[8]_i_1_n_11 ,\total_bytes_recved_reg[8]_i_1_n_12 ,\total_bytes_recved_reg[8]_i_1_n_13 ,\total_bytes_recved_reg[8]_i_1_n_14 ,\total_bytes_recved_reg[8]_i_1_n_15 }),
        .S(total_bytes_recved_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_recved_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[18]),
        .CLR(rst_i),
        .D(\total_bytes_recved_reg[8]_i_1_n_14 ),
        .Q(total_bytes_recved_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \total_bytes_transed[0]_i_2 
       (.I0(total_bytes_transed_reg[0]),
        .O(\total_bytes_transed[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[0]_i_1_n_0 ,\total_bytes_transed_reg[0]_i_1_n_1 ,\total_bytes_transed_reg[0]_i_1_n_2 ,\total_bytes_transed_reg[0]_i_1_n_3 ,\total_bytes_transed_reg[0]_i_1_n_4 ,\total_bytes_transed_reg[0]_i_1_n_5 ,\total_bytes_transed_reg[0]_i_1_n_6 ,\total_bytes_transed_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\total_bytes_transed_reg[0]_i_1_n_8 ,\total_bytes_transed_reg[0]_i_1_n_9 ,\total_bytes_transed_reg[0]_i_1_n_10 ,\total_bytes_transed_reg[0]_i_1_n_11 ,\total_bytes_transed_reg[0]_i_1_n_12 ,\total_bytes_transed_reg[0]_i_1_n_13 ,\total_bytes_transed_reg[0]_i_1_n_14 ,\total_bytes_transed_reg[0]_i_1_n_15 }),
        .S({total_bytes_transed_reg[7:1],\total_bytes_transed[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[16]_i_1 
       (.CI(\total_bytes_transed_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[16]_i_1_n_0 ,\total_bytes_transed_reg[16]_i_1_n_1 ,\total_bytes_transed_reg[16]_i_1_n_2 ,\total_bytes_transed_reg[16]_i_1_n_3 ,\total_bytes_transed_reg[16]_i_1_n_4 ,\total_bytes_transed_reg[16]_i_1_n_5 ,\total_bytes_transed_reg[16]_i_1_n_6 ,\total_bytes_transed_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[16]_i_1_n_8 ,\total_bytes_transed_reg[16]_i_1_n_9 ,\total_bytes_transed_reg[16]_i_1_n_10 ,\total_bytes_transed_reg[16]_i_1_n_11 ,\total_bytes_transed_reg[16]_i_1_n_12 ,\total_bytes_transed_reg[16]_i_1_n_13 ,\total_bytes_transed_reg[16]_i_1_n_14 ,\total_bytes_transed_reg[16]_i_1_n_15 }),
        .S(total_bytes_transed_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[16]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[24]_i_1 
       (.CI(\total_bytes_transed_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[24]_i_1_n_0 ,\total_bytes_transed_reg[24]_i_1_n_1 ,\total_bytes_transed_reg[24]_i_1_n_2 ,\total_bytes_transed_reg[24]_i_1_n_3 ,\total_bytes_transed_reg[24]_i_1_n_4 ,\total_bytes_transed_reg[24]_i_1_n_5 ,\total_bytes_transed_reg[24]_i_1_n_6 ,\total_bytes_transed_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[24]_i_1_n_8 ,\total_bytes_transed_reg[24]_i_1_n_9 ,\total_bytes_transed_reg[24]_i_1_n_10 ,\total_bytes_transed_reg[24]_i_1_n_11 ,\total_bytes_transed_reg[24]_i_1_n_12 ,\total_bytes_transed_reg[24]_i_1_n_13 ,\total_bytes_transed_reg[24]_i_1_n_14 ,\total_bytes_transed_reg[24]_i_1_n_15 }),
        .S(total_bytes_transed_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[24]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[32]_i_1 
       (.CI(\total_bytes_transed_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[32]_i_1_n_0 ,\total_bytes_transed_reg[32]_i_1_n_1 ,\total_bytes_transed_reg[32]_i_1_n_2 ,\total_bytes_transed_reg[32]_i_1_n_3 ,\total_bytes_transed_reg[32]_i_1_n_4 ,\total_bytes_transed_reg[32]_i_1_n_5 ,\total_bytes_transed_reg[32]_i_1_n_6 ,\total_bytes_transed_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[32]_i_1_n_8 ,\total_bytes_transed_reg[32]_i_1_n_9 ,\total_bytes_transed_reg[32]_i_1_n_10 ,\total_bytes_transed_reg[32]_i_1_n_11 ,\total_bytes_transed_reg[32]_i_1_n_12 ,\total_bytes_transed_reg[32]_i_1_n_13 ,\total_bytes_transed_reg[32]_i_1_n_14 ,\total_bytes_transed_reg[32]_i_1_n_15 }),
        .S(total_bytes_transed_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[32]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[40]_i_1 
       (.CI(\total_bytes_transed_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[40]_i_1_n_0 ,\total_bytes_transed_reg[40]_i_1_n_1 ,\total_bytes_transed_reg[40]_i_1_n_2 ,\total_bytes_transed_reg[40]_i_1_n_3 ,\total_bytes_transed_reg[40]_i_1_n_4 ,\total_bytes_transed_reg[40]_i_1_n_5 ,\total_bytes_transed_reg[40]_i_1_n_6 ,\total_bytes_transed_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[40]_i_1_n_8 ,\total_bytes_transed_reg[40]_i_1_n_9 ,\total_bytes_transed_reg[40]_i_1_n_10 ,\total_bytes_transed_reg[40]_i_1_n_11 ,\total_bytes_transed_reg[40]_i_1_n_12 ,\total_bytes_transed_reg[40]_i_1_n_13 ,\total_bytes_transed_reg[40]_i_1_n_14 ,\total_bytes_transed_reg[40]_i_1_n_15 }),
        .S(total_bytes_transed_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[40]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[48]_i_1 
       (.CI(\total_bytes_transed_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[48]_i_1_n_0 ,\total_bytes_transed_reg[48]_i_1_n_1 ,\total_bytes_transed_reg[48]_i_1_n_2 ,\total_bytes_transed_reg[48]_i_1_n_3 ,\total_bytes_transed_reg[48]_i_1_n_4 ,\total_bytes_transed_reg[48]_i_1_n_5 ,\total_bytes_transed_reg[48]_i_1_n_6 ,\total_bytes_transed_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[48]_i_1_n_8 ,\total_bytes_transed_reg[48]_i_1_n_9 ,\total_bytes_transed_reg[48]_i_1_n_10 ,\total_bytes_transed_reg[48]_i_1_n_11 ,\total_bytes_transed_reg[48]_i_1_n_12 ,\total_bytes_transed_reg[48]_i_1_n_13 ,\total_bytes_transed_reg[48]_i_1_n_14 ,\total_bytes_transed_reg[48]_i_1_n_15 }),
        .S(total_bytes_transed_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[48]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[56]_i_1 
       (.CI(\total_bytes_transed_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_total_bytes_transed_reg[56]_i_1_CO_UNCONNECTED [7],\total_bytes_transed_reg[56]_i_1_n_1 ,\total_bytes_transed_reg[56]_i_1_n_2 ,\total_bytes_transed_reg[56]_i_1_n_3 ,\total_bytes_transed_reg[56]_i_1_n_4 ,\total_bytes_transed_reg[56]_i_1_n_5 ,\total_bytes_transed_reg[56]_i_1_n_6 ,\total_bytes_transed_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[56]_i_1_n_8 ,\total_bytes_transed_reg[56]_i_1_n_9 ,\total_bytes_transed_reg[56]_i_1_n_10 ,\total_bytes_transed_reg[56]_i_1_n_11 ,\total_bytes_transed_reg[56]_i_1_n_12 ,\total_bytes_transed_reg[56]_i_1_n_13 ,\total_bytes_transed_reg[56]_i_1_n_14 ,\total_bytes_transed_reg[56]_i_1_n_15 }),
        .S(total_bytes_transed_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_13 ),
        .Q(total_bytes_transed_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_12 ),
        .Q(total_bytes_transed_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_11 ),
        .Q(total_bytes_transed_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_10 ),
        .Q(total_bytes_transed_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[56]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_9 ),
        .Q(total_bytes_transed_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[0]_i_1_n_8 ),
        .Q(total_bytes_transed_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_15 ),
        .Q(total_bytes_transed_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \total_bytes_transed_reg[8]_i_1 
       (.CI(\total_bytes_transed_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\total_bytes_transed_reg[8]_i_1_n_0 ,\total_bytes_transed_reg[8]_i_1_n_1 ,\total_bytes_transed_reg[8]_i_1_n_2 ,\total_bytes_transed_reg[8]_i_1_n_3 ,\total_bytes_transed_reg[8]_i_1_n_4 ,\total_bytes_transed_reg[8]_i_1_n_5 ,\total_bytes_transed_reg[8]_i_1_n_6 ,\total_bytes_transed_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\total_bytes_transed_reg[8]_i_1_n_8 ,\total_bytes_transed_reg[8]_i_1_n_9 ,\total_bytes_transed_reg[8]_i_1_n_10 ,\total_bytes_transed_reg[8]_i_1_n_11 ,\total_bytes_transed_reg[8]_i_1_n_12 ,\total_bytes_transed_reg[8]_i_1_n_13 ,\total_bytes_transed_reg[8]_i_1_n_14 ,\total_bytes_transed_reg[8]_i_1_n_15 }),
        .S(total_bytes_transed_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \total_bytes_transed_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[0]),
        .CLR(rst_i),
        .D(\total_bytes_transed_reg[8]_i_1_n_14 ),
        .Q(total_bytes_transed_reg[9]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \trans_config[31]_i_1 
       (.I0(\recv_config0_reg[0]_0 ),
        .I1(out[9]),
        .I2(\stat_rd_data_reg[63]_1 ),
        .I3(\trans_config[31]_i_2_n_0 ),
        .I4(\recv_config1[31]_i_4_n_0 ),
        .I5(out[7]),
        .O(\trans_config[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \trans_config[31]_i_2 
       (.I0(out[8]),
        .I1(out[0]),
        .I2(out[5]),
        .I3(out[6]),
        .O(\trans_config[31]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[0] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[0]),
        .Q(\trans_config_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[10] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[10]),
        .Q(\trans_config_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[11] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[11]),
        .Q(\trans_config_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[12] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[12]),
        .Q(\trans_config_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[13] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[13]),
        .Q(\trans_config_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[14] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[14]),
        .Q(\trans_config_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[15] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[15]),
        .Q(\trans_config_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[16] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[16]),
        .Q(\trans_config_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[17] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[17]),
        .Q(\trans_config_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[18] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[18]),
        .Q(\trans_config_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[19] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[19]),
        .Q(\trans_config_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[1] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[1]),
        .Q(\trans_config_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[20] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[20]),
        .Q(\trans_config_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[21] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[21]),
        .Q(\trans_config_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[22] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[22]),
        .Q(\trans_config_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[23] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[23]),
        .Q(\trans_config_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[24] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[24]),
        .Q(cfgTxRegData[1]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[25] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[25]),
        .Q(cfgTxRegData[2]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[26] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[26]),
        .Q(cfgTxRegData[3]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[27] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[27]),
        .Q(cfgTxRegData[4]));
  FDPE #(
    .INIT(1'b1)) 
    \trans_config_reg[28] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .D(mgmt_wr_data[28]),
        .PRE(rst_i),
        .Q(cfgTxRegData[5]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[29] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[29]),
        .Q(cfgTxRegData[6]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[2] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[2]),
        .Q(\trans_config_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[30] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[30]),
        .Q(cfgTxRegData[7]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[31] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[31]),
        .Q(cfgTxRegData[8]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[3] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[3]),
        .Q(\trans_config_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[4] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[4]),
        .Q(\trans_config_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[5] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[5]),
        .Q(\trans_config_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[6] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[6]),
        .Q(\trans_config_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[7] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[7]),
        .Q(\trans_config_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[8] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[8]),
        .Q(\trans_config_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_config_reg[9] 
       (.C(clk_i),
        .CE(\trans_config[31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(mgmt_wr_data[9]),
        .Q(\trans_config_reg_n_0_[9] ));
  LUT1 #(
    .INIT(2'h1)) 
    \underrun_error[0]_i_2 
       (.I0(underrun_error_reg[0]),
        .O(\underrun_error[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[0] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_15 ),
        .Q(underrun_error_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[0]_i_1_n_0 ,\underrun_error_reg[0]_i_1_n_1 ,\underrun_error_reg[0]_i_1_n_2 ,\underrun_error_reg[0]_i_1_n_3 ,\underrun_error_reg[0]_i_1_n_4 ,\underrun_error_reg[0]_i_1_n_5 ,\underrun_error_reg[0]_i_1_n_6 ,\underrun_error_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\underrun_error_reg[0]_i_1_n_8 ,\underrun_error_reg[0]_i_1_n_9 ,\underrun_error_reg[0]_i_1_n_10 ,\underrun_error_reg[0]_i_1_n_11 ,\underrun_error_reg[0]_i_1_n_12 ,\underrun_error_reg[0]_i_1_n_13 ,\underrun_error_reg[0]_i_1_n_14 ,\underrun_error_reg[0]_i_1_n_15 }),
        .S({underrun_error_reg[7:1],\underrun_error[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[10] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_13 ),
        .Q(underrun_error_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[11] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_12 ),
        .Q(underrun_error_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[12] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_11 ),
        .Q(underrun_error_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[13] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_10 ),
        .Q(underrun_error_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[14] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_9 ),
        .Q(underrun_error_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[15] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_8 ),
        .Q(underrun_error_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[16] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_15 ),
        .Q(underrun_error_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[16]_i_1 
       (.CI(\underrun_error_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[16]_i_1_n_0 ,\underrun_error_reg[16]_i_1_n_1 ,\underrun_error_reg[16]_i_1_n_2 ,\underrun_error_reg[16]_i_1_n_3 ,\underrun_error_reg[16]_i_1_n_4 ,\underrun_error_reg[16]_i_1_n_5 ,\underrun_error_reg[16]_i_1_n_6 ,\underrun_error_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[16]_i_1_n_8 ,\underrun_error_reg[16]_i_1_n_9 ,\underrun_error_reg[16]_i_1_n_10 ,\underrun_error_reg[16]_i_1_n_11 ,\underrun_error_reg[16]_i_1_n_12 ,\underrun_error_reg[16]_i_1_n_13 ,\underrun_error_reg[16]_i_1_n_14 ,\underrun_error_reg[16]_i_1_n_15 }),
        .S(underrun_error_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[17] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_14 ),
        .Q(underrun_error_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[18] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_13 ),
        .Q(underrun_error_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[19] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_12 ),
        .Q(underrun_error_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[1] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_14 ),
        .Q(underrun_error_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[20] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_11 ),
        .Q(underrun_error_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[21] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_10 ),
        .Q(underrun_error_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[22] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_9 ),
        .Q(underrun_error_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[23] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[16]_i_1_n_8 ),
        .Q(underrun_error_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[24] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_15 ),
        .Q(underrun_error_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[24]_i_1 
       (.CI(\underrun_error_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[24]_i_1_n_0 ,\underrun_error_reg[24]_i_1_n_1 ,\underrun_error_reg[24]_i_1_n_2 ,\underrun_error_reg[24]_i_1_n_3 ,\underrun_error_reg[24]_i_1_n_4 ,\underrun_error_reg[24]_i_1_n_5 ,\underrun_error_reg[24]_i_1_n_6 ,\underrun_error_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[24]_i_1_n_8 ,\underrun_error_reg[24]_i_1_n_9 ,\underrun_error_reg[24]_i_1_n_10 ,\underrun_error_reg[24]_i_1_n_11 ,\underrun_error_reg[24]_i_1_n_12 ,\underrun_error_reg[24]_i_1_n_13 ,\underrun_error_reg[24]_i_1_n_14 ,\underrun_error_reg[24]_i_1_n_15 }),
        .S(underrun_error_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[25] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_14 ),
        .Q(underrun_error_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[26] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_13 ),
        .Q(underrun_error_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[27] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_12 ),
        .Q(underrun_error_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[28] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_11 ),
        .Q(underrun_error_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[29] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_10 ),
        .Q(underrun_error_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[2] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_13 ),
        .Q(underrun_error_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[30] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_9 ),
        .Q(underrun_error_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[31] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[24]_i_1_n_8 ),
        .Q(underrun_error_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[32] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_15 ),
        .Q(underrun_error_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[32]_i_1 
       (.CI(\underrun_error_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[32]_i_1_n_0 ,\underrun_error_reg[32]_i_1_n_1 ,\underrun_error_reg[32]_i_1_n_2 ,\underrun_error_reg[32]_i_1_n_3 ,\underrun_error_reg[32]_i_1_n_4 ,\underrun_error_reg[32]_i_1_n_5 ,\underrun_error_reg[32]_i_1_n_6 ,\underrun_error_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[32]_i_1_n_8 ,\underrun_error_reg[32]_i_1_n_9 ,\underrun_error_reg[32]_i_1_n_10 ,\underrun_error_reg[32]_i_1_n_11 ,\underrun_error_reg[32]_i_1_n_12 ,\underrun_error_reg[32]_i_1_n_13 ,\underrun_error_reg[32]_i_1_n_14 ,\underrun_error_reg[32]_i_1_n_15 }),
        .S(underrun_error_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[33] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_14 ),
        .Q(underrun_error_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[34] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_13 ),
        .Q(underrun_error_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[35] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_12 ),
        .Q(underrun_error_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[36] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_11 ),
        .Q(underrun_error_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[37] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_10 ),
        .Q(underrun_error_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[38] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_9 ),
        .Q(underrun_error_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[39] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[32]_i_1_n_8 ),
        .Q(underrun_error_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[3] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_12 ),
        .Q(underrun_error_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[40] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_15 ),
        .Q(underrun_error_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[40]_i_1 
       (.CI(\underrun_error_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[40]_i_1_n_0 ,\underrun_error_reg[40]_i_1_n_1 ,\underrun_error_reg[40]_i_1_n_2 ,\underrun_error_reg[40]_i_1_n_3 ,\underrun_error_reg[40]_i_1_n_4 ,\underrun_error_reg[40]_i_1_n_5 ,\underrun_error_reg[40]_i_1_n_6 ,\underrun_error_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[40]_i_1_n_8 ,\underrun_error_reg[40]_i_1_n_9 ,\underrun_error_reg[40]_i_1_n_10 ,\underrun_error_reg[40]_i_1_n_11 ,\underrun_error_reg[40]_i_1_n_12 ,\underrun_error_reg[40]_i_1_n_13 ,\underrun_error_reg[40]_i_1_n_14 ,\underrun_error_reg[40]_i_1_n_15 }),
        .S(underrun_error_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[41] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_14 ),
        .Q(underrun_error_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[42] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_13 ),
        .Q(underrun_error_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[43] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_12 ),
        .Q(underrun_error_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[44] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_11 ),
        .Q(underrun_error_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[45] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_10 ),
        .Q(underrun_error_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[46] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_9 ),
        .Q(underrun_error_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[47] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[40]_i_1_n_8 ),
        .Q(underrun_error_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[48] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_15 ),
        .Q(underrun_error_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[48]_i_1 
       (.CI(\underrun_error_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[48]_i_1_n_0 ,\underrun_error_reg[48]_i_1_n_1 ,\underrun_error_reg[48]_i_1_n_2 ,\underrun_error_reg[48]_i_1_n_3 ,\underrun_error_reg[48]_i_1_n_4 ,\underrun_error_reg[48]_i_1_n_5 ,\underrun_error_reg[48]_i_1_n_6 ,\underrun_error_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[48]_i_1_n_8 ,\underrun_error_reg[48]_i_1_n_9 ,\underrun_error_reg[48]_i_1_n_10 ,\underrun_error_reg[48]_i_1_n_11 ,\underrun_error_reg[48]_i_1_n_12 ,\underrun_error_reg[48]_i_1_n_13 ,\underrun_error_reg[48]_i_1_n_14 ,\underrun_error_reg[48]_i_1_n_15 }),
        .S(underrun_error_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[49] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_14 ),
        .Q(underrun_error_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[4] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_11 ),
        .Q(underrun_error_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[50] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_13 ),
        .Q(underrun_error_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[51] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_12 ),
        .Q(underrun_error_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[52] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_11 ),
        .Q(underrun_error_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[53] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_10 ),
        .Q(underrun_error_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[54] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_9 ),
        .Q(underrun_error_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[55] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[48]_i_1_n_8 ),
        .Q(underrun_error_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[56] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_15 ),
        .Q(underrun_error_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[56]_i_1 
       (.CI(\underrun_error_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_underrun_error_reg[56]_i_1_CO_UNCONNECTED [7],\underrun_error_reg[56]_i_1_n_1 ,\underrun_error_reg[56]_i_1_n_2 ,\underrun_error_reg[56]_i_1_n_3 ,\underrun_error_reg[56]_i_1_n_4 ,\underrun_error_reg[56]_i_1_n_5 ,\underrun_error_reg[56]_i_1_n_6 ,\underrun_error_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[56]_i_1_n_8 ,\underrun_error_reg[56]_i_1_n_9 ,\underrun_error_reg[56]_i_1_n_10 ,\underrun_error_reg[56]_i_1_n_11 ,\underrun_error_reg[56]_i_1_n_12 ,\underrun_error_reg[56]_i_1_n_13 ,\underrun_error_reg[56]_i_1_n_14 ,\underrun_error_reg[56]_i_1_n_15 }),
        .S(underrun_error_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[57] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_14 ),
        .Q(underrun_error_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[58] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_13 ),
        .Q(underrun_error_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[59] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_12 ),
        .Q(underrun_error_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[5] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_10 ),
        .Q(underrun_error_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[60] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_11 ),
        .Q(underrun_error_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[61] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_10 ),
        .Q(underrun_error_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[62] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_9 ),
        .Q(underrun_error_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[63] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[56]_i_1_n_8 ),
        .Q(underrun_error_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[6] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_9 ),
        .Q(underrun_error_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[7] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[0]_i_1_n_8 ),
        .Q(underrun_error_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[8] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_15 ),
        .Q(underrun_error_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \underrun_error_reg[8]_i_1 
       (.CI(\underrun_error_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\underrun_error_reg[8]_i_1_n_0 ,\underrun_error_reg[8]_i_1_n_1 ,\underrun_error_reg[8]_i_1_n_2 ,\underrun_error_reg[8]_i_1_n_3 ,\underrun_error_reg[8]_i_1_n_4 ,\underrun_error_reg[8]_i_1_n_5 ,\underrun_error_reg[8]_i_1_n_6 ,\underrun_error_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\underrun_error_reg[8]_i_1_n_8 ,\underrun_error_reg[8]_i_1_n_9 ,\underrun_error_reg[8]_i_1_n_10 ,\underrun_error_reg[8]_i_1_n_11 ,\underrun_error_reg[8]_i_1_n_12 ,\underrun_error_reg[8]_i_1_n_13 ,\underrun_error_reg[8]_i_1_n_14 ,\underrun_error_reg[8]_i_1_n_15 }),
        .S(underrun_error_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \underrun_error_reg[9] 
       (.C(clk_i),
        .CE(txStatRegPlus[4]),
        .CLR(rst_i),
        .D(\underrun_error_reg[8]_i_1_n_14 ),
        .Q(underrun_error_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \undersize_frame[0]_i_2 
       (.I0(undersize_frame_reg[0]),
        .O(\undersize_frame[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_15 ),
        .Q(undersize_frame_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[0]_i_1_n_0 ,\undersize_frame_reg[0]_i_1_n_1 ,\undersize_frame_reg[0]_i_1_n_2 ,\undersize_frame_reg[0]_i_1_n_3 ,\undersize_frame_reg[0]_i_1_n_4 ,\undersize_frame_reg[0]_i_1_n_5 ,\undersize_frame_reg[0]_i_1_n_6 ,\undersize_frame_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\undersize_frame_reg[0]_i_1_n_8 ,\undersize_frame_reg[0]_i_1_n_9 ,\undersize_frame_reg[0]_i_1_n_10 ,\undersize_frame_reg[0]_i_1_n_11 ,\undersize_frame_reg[0]_i_1_n_12 ,\undersize_frame_reg[0]_i_1_n_13 ,\undersize_frame_reg[0]_i_1_n_14 ,\undersize_frame_reg[0]_i_1_n_15 }),
        .S({undersize_frame_reg[7:1],\undersize_frame[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_13 ),
        .Q(undersize_frame_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_12 ),
        .Q(undersize_frame_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_11 ),
        .Q(undersize_frame_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_10 ),
        .Q(undersize_frame_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_9 ),
        .Q(undersize_frame_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_8 ),
        .Q(undersize_frame_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_15 ),
        .Q(undersize_frame_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[16]_i_1 
       (.CI(\undersize_frame_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[16]_i_1_n_0 ,\undersize_frame_reg[16]_i_1_n_1 ,\undersize_frame_reg[16]_i_1_n_2 ,\undersize_frame_reg[16]_i_1_n_3 ,\undersize_frame_reg[16]_i_1_n_4 ,\undersize_frame_reg[16]_i_1_n_5 ,\undersize_frame_reg[16]_i_1_n_6 ,\undersize_frame_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[16]_i_1_n_8 ,\undersize_frame_reg[16]_i_1_n_9 ,\undersize_frame_reg[16]_i_1_n_10 ,\undersize_frame_reg[16]_i_1_n_11 ,\undersize_frame_reg[16]_i_1_n_12 ,\undersize_frame_reg[16]_i_1_n_13 ,\undersize_frame_reg[16]_i_1_n_14 ,\undersize_frame_reg[16]_i_1_n_15 }),
        .S(undersize_frame_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_14 ),
        .Q(undersize_frame_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_13 ),
        .Q(undersize_frame_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_12 ),
        .Q(undersize_frame_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_14 ),
        .Q(undersize_frame_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_11 ),
        .Q(undersize_frame_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_10 ),
        .Q(undersize_frame_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_9 ),
        .Q(undersize_frame_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[16]_i_1_n_8 ),
        .Q(undersize_frame_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_15 ),
        .Q(undersize_frame_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[24]_i_1 
       (.CI(\undersize_frame_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[24]_i_1_n_0 ,\undersize_frame_reg[24]_i_1_n_1 ,\undersize_frame_reg[24]_i_1_n_2 ,\undersize_frame_reg[24]_i_1_n_3 ,\undersize_frame_reg[24]_i_1_n_4 ,\undersize_frame_reg[24]_i_1_n_5 ,\undersize_frame_reg[24]_i_1_n_6 ,\undersize_frame_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[24]_i_1_n_8 ,\undersize_frame_reg[24]_i_1_n_9 ,\undersize_frame_reg[24]_i_1_n_10 ,\undersize_frame_reg[24]_i_1_n_11 ,\undersize_frame_reg[24]_i_1_n_12 ,\undersize_frame_reg[24]_i_1_n_13 ,\undersize_frame_reg[24]_i_1_n_14 ,\undersize_frame_reg[24]_i_1_n_15 }),
        .S(undersize_frame_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_14 ),
        .Q(undersize_frame_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_13 ),
        .Q(undersize_frame_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_12 ),
        .Q(undersize_frame_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_11 ),
        .Q(undersize_frame_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_10 ),
        .Q(undersize_frame_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_13 ),
        .Q(undersize_frame_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_9 ),
        .Q(undersize_frame_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[24]_i_1_n_8 ),
        .Q(undersize_frame_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_15 ),
        .Q(undersize_frame_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[32]_i_1 
       (.CI(\undersize_frame_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[32]_i_1_n_0 ,\undersize_frame_reg[32]_i_1_n_1 ,\undersize_frame_reg[32]_i_1_n_2 ,\undersize_frame_reg[32]_i_1_n_3 ,\undersize_frame_reg[32]_i_1_n_4 ,\undersize_frame_reg[32]_i_1_n_5 ,\undersize_frame_reg[32]_i_1_n_6 ,\undersize_frame_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[32]_i_1_n_8 ,\undersize_frame_reg[32]_i_1_n_9 ,\undersize_frame_reg[32]_i_1_n_10 ,\undersize_frame_reg[32]_i_1_n_11 ,\undersize_frame_reg[32]_i_1_n_12 ,\undersize_frame_reg[32]_i_1_n_13 ,\undersize_frame_reg[32]_i_1_n_14 ,\undersize_frame_reg[32]_i_1_n_15 }),
        .S(undersize_frame_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_14 ),
        .Q(undersize_frame_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_13 ),
        .Q(undersize_frame_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_12 ),
        .Q(undersize_frame_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_11 ),
        .Q(undersize_frame_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_10 ),
        .Q(undersize_frame_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_9 ),
        .Q(undersize_frame_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[32]_i_1_n_8 ),
        .Q(undersize_frame_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_12 ),
        .Q(undersize_frame_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_15 ),
        .Q(undersize_frame_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[40]_i_1 
       (.CI(\undersize_frame_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[40]_i_1_n_0 ,\undersize_frame_reg[40]_i_1_n_1 ,\undersize_frame_reg[40]_i_1_n_2 ,\undersize_frame_reg[40]_i_1_n_3 ,\undersize_frame_reg[40]_i_1_n_4 ,\undersize_frame_reg[40]_i_1_n_5 ,\undersize_frame_reg[40]_i_1_n_6 ,\undersize_frame_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[40]_i_1_n_8 ,\undersize_frame_reg[40]_i_1_n_9 ,\undersize_frame_reg[40]_i_1_n_10 ,\undersize_frame_reg[40]_i_1_n_11 ,\undersize_frame_reg[40]_i_1_n_12 ,\undersize_frame_reg[40]_i_1_n_13 ,\undersize_frame_reg[40]_i_1_n_14 ,\undersize_frame_reg[40]_i_1_n_15 }),
        .S(undersize_frame_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_14 ),
        .Q(undersize_frame_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_13 ),
        .Q(undersize_frame_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_12 ),
        .Q(undersize_frame_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_11 ),
        .Q(undersize_frame_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_10 ),
        .Q(undersize_frame_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_9 ),
        .Q(undersize_frame_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[40]_i_1_n_8 ),
        .Q(undersize_frame_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_15 ),
        .Q(undersize_frame_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[48]_i_1 
       (.CI(\undersize_frame_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[48]_i_1_n_0 ,\undersize_frame_reg[48]_i_1_n_1 ,\undersize_frame_reg[48]_i_1_n_2 ,\undersize_frame_reg[48]_i_1_n_3 ,\undersize_frame_reg[48]_i_1_n_4 ,\undersize_frame_reg[48]_i_1_n_5 ,\undersize_frame_reg[48]_i_1_n_6 ,\undersize_frame_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[48]_i_1_n_8 ,\undersize_frame_reg[48]_i_1_n_9 ,\undersize_frame_reg[48]_i_1_n_10 ,\undersize_frame_reg[48]_i_1_n_11 ,\undersize_frame_reg[48]_i_1_n_12 ,\undersize_frame_reg[48]_i_1_n_13 ,\undersize_frame_reg[48]_i_1_n_14 ,\undersize_frame_reg[48]_i_1_n_15 }),
        .S(undersize_frame_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_14 ),
        .Q(undersize_frame_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_11 ),
        .Q(undersize_frame_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_13 ),
        .Q(undersize_frame_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_12 ),
        .Q(undersize_frame_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_11 ),
        .Q(undersize_frame_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_10 ),
        .Q(undersize_frame_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_9 ),
        .Q(undersize_frame_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[48]_i_1_n_8 ),
        .Q(undersize_frame_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_15 ),
        .Q(undersize_frame_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[56]_i_1 
       (.CI(\undersize_frame_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_undersize_frame_reg[56]_i_1_CO_UNCONNECTED [7],\undersize_frame_reg[56]_i_1_n_1 ,\undersize_frame_reg[56]_i_1_n_2 ,\undersize_frame_reg[56]_i_1_n_3 ,\undersize_frame_reg[56]_i_1_n_4 ,\undersize_frame_reg[56]_i_1_n_5 ,\undersize_frame_reg[56]_i_1_n_6 ,\undersize_frame_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[56]_i_1_n_8 ,\undersize_frame_reg[56]_i_1_n_9 ,\undersize_frame_reg[56]_i_1_n_10 ,\undersize_frame_reg[56]_i_1_n_11 ,\undersize_frame_reg[56]_i_1_n_12 ,\undersize_frame_reg[56]_i_1_n_13 ,\undersize_frame_reg[56]_i_1_n_14 ,\undersize_frame_reg[56]_i_1_n_15 }),
        .S(undersize_frame_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_14 ),
        .Q(undersize_frame_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_13 ),
        .Q(undersize_frame_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_12 ),
        .Q(undersize_frame_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_10 ),
        .Q(undersize_frame_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_11 ),
        .Q(undersize_frame_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_10 ),
        .Q(undersize_frame_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_9 ),
        .Q(undersize_frame_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[56]_i_1_n_8 ),
        .Q(undersize_frame_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_9 ),
        .Q(undersize_frame_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[0]_i_1_n_8 ),
        .Q(undersize_frame_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_15 ),
        .Q(undersize_frame_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \undersize_frame_reg[8]_i_1 
       (.CI(\undersize_frame_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\undersize_frame_reg[8]_i_1_n_0 ,\undersize_frame_reg[8]_i_1_n_1 ,\undersize_frame_reg[8]_i_1_n_2 ,\undersize_frame_reg[8]_i_1_n_3 ,\undersize_frame_reg[8]_i_1_n_4 ,\undersize_frame_reg[8]_i_1_n_5 ,\undersize_frame_reg[8]_i_1_n_6 ,\undersize_frame_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\undersize_frame_reg[8]_i_1_n_8 ,\undersize_frame_reg[8]_i_1_n_9 ,\undersize_frame_reg[8]_i_1_n_10 ,\undersize_frame_reg[8]_i_1_n_11 ,\undersize_frame_reg[8]_i_1_n_12 ,\undersize_frame_reg[8]_i_1_n_13 ,\undersize_frame_reg[8]_i_1_n_14 ,\undersize_frame_reg[8]_i_1_n_15 }),
        .S(undersize_frame_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \undersize_frame_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[16]),
        .CLR(rst_i),
        .D(\undersize_frame_reg[8]_i_1_n_14 ),
        .Q(undersize_frame_reg[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \unsupported_control_frame[0]_i_2 
       (.I0(unsupported_control_frame_reg[0]),
        .O(\unsupported_control_frame[0]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[0] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[0]_i_1_n_0 ,\unsupported_control_frame_reg[0]_i_1_n_1 ,\unsupported_control_frame_reg[0]_i_1_n_2 ,\unsupported_control_frame_reg[0]_i_1_n_3 ,\unsupported_control_frame_reg[0]_i_1_n_4 ,\unsupported_control_frame_reg[0]_i_1_n_5 ,\unsupported_control_frame_reg[0]_i_1_n_6 ,\unsupported_control_frame_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}),
        .O({\unsupported_control_frame_reg[0]_i_1_n_8 ,\unsupported_control_frame_reg[0]_i_1_n_9 ,\unsupported_control_frame_reg[0]_i_1_n_10 ,\unsupported_control_frame_reg[0]_i_1_n_11 ,\unsupported_control_frame_reg[0]_i_1_n_12 ,\unsupported_control_frame_reg[0]_i_1_n_13 ,\unsupported_control_frame_reg[0]_i_1_n_14 ,\unsupported_control_frame_reg[0]_i_1_n_15 }),
        .S({unsupported_control_frame_reg[7:1],\unsupported_control_frame[0]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[10] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[11] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[12] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[13] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[14] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[15] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[16] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[16]_i_1 
       (.CI(\unsupported_control_frame_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[16]_i_1_n_0 ,\unsupported_control_frame_reg[16]_i_1_n_1 ,\unsupported_control_frame_reg[16]_i_1_n_2 ,\unsupported_control_frame_reg[16]_i_1_n_3 ,\unsupported_control_frame_reg[16]_i_1_n_4 ,\unsupported_control_frame_reg[16]_i_1_n_5 ,\unsupported_control_frame_reg[16]_i_1_n_6 ,\unsupported_control_frame_reg[16]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[16]_i_1_n_8 ,\unsupported_control_frame_reg[16]_i_1_n_9 ,\unsupported_control_frame_reg[16]_i_1_n_10 ,\unsupported_control_frame_reg[16]_i_1_n_11 ,\unsupported_control_frame_reg[16]_i_1_n_12 ,\unsupported_control_frame_reg[16]_i_1_n_13 ,\unsupported_control_frame_reg[16]_i_1_n_14 ,\unsupported_control_frame_reg[16]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[23:16]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[17] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[18] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[19] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[1] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[20] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[21] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[22] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[23] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[16]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[24] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[24]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[24]_i_1 
       (.CI(\unsupported_control_frame_reg[16]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[24]_i_1_n_0 ,\unsupported_control_frame_reg[24]_i_1_n_1 ,\unsupported_control_frame_reg[24]_i_1_n_2 ,\unsupported_control_frame_reg[24]_i_1_n_3 ,\unsupported_control_frame_reg[24]_i_1_n_4 ,\unsupported_control_frame_reg[24]_i_1_n_5 ,\unsupported_control_frame_reg[24]_i_1_n_6 ,\unsupported_control_frame_reg[24]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[24]_i_1_n_8 ,\unsupported_control_frame_reg[24]_i_1_n_9 ,\unsupported_control_frame_reg[24]_i_1_n_10 ,\unsupported_control_frame_reg[24]_i_1_n_11 ,\unsupported_control_frame_reg[24]_i_1_n_12 ,\unsupported_control_frame_reg[24]_i_1_n_13 ,\unsupported_control_frame_reg[24]_i_1_n_14 ,\unsupported_control_frame_reg[24]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[31:24]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[25] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[26] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[27] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[28] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[29] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[2] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[30] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[31] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[24]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[32] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[32]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[32]_i_1 
       (.CI(\unsupported_control_frame_reg[24]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[32]_i_1_n_0 ,\unsupported_control_frame_reg[32]_i_1_n_1 ,\unsupported_control_frame_reg[32]_i_1_n_2 ,\unsupported_control_frame_reg[32]_i_1_n_3 ,\unsupported_control_frame_reg[32]_i_1_n_4 ,\unsupported_control_frame_reg[32]_i_1_n_5 ,\unsupported_control_frame_reg[32]_i_1_n_6 ,\unsupported_control_frame_reg[32]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[32]_i_1_n_8 ,\unsupported_control_frame_reg[32]_i_1_n_9 ,\unsupported_control_frame_reg[32]_i_1_n_10 ,\unsupported_control_frame_reg[32]_i_1_n_11 ,\unsupported_control_frame_reg[32]_i_1_n_12 ,\unsupported_control_frame_reg[32]_i_1_n_13 ,\unsupported_control_frame_reg[32]_i_1_n_14 ,\unsupported_control_frame_reg[32]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[39:32]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[33] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[34] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[35] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[36] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[37] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[38] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[39] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[32]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[3] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[40] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[40]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[40]_i_1 
       (.CI(\unsupported_control_frame_reg[32]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[40]_i_1_n_0 ,\unsupported_control_frame_reg[40]_i_1_n_1 ,\unsupported_control_frame_reg[40]_i_1_n_2 ,\unsupported_control_frame_reg[40]_i_1_n_3 ,\unsupported_control_frame_reg[40]_i_1_n_4 ,\unsupported_control_frame_reg[40]_i_1_n_5 ,\unsupported_control_frame_reg[40]_i_1_n_6 ,\unsupported_control_frame_reg[40]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[40]_i_1_n_8 ,\unsupported_control_frame_reg[40]_i_1_n_9 ,\unsupported_control_frame_reg[40]_i_1_n_10 ,\unsupported_control_frame_reg[40]_i_1_n_11 ,\unsupported_control_frame_reg[40]_i_1_n_12 ,\unsupported_control_frame_reg[40]_i_1_n_13 ,\unsupported_control_frame_reg[40]_i_1_n_14 ,\unsupported_control_frame_reg[40]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[47:40]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[41] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[42] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[43] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[44] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[45] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[46] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[47] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[40]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[48] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[48]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[48]_i_1 
       (.CI(\unsupported_control_frame_reg[40]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[48]_i_1_n_0 ,\unsupported_control_frame_reg[48]_i_1_n_1 ,\unsupported_control_frame_reg[48]_i_1_n_2 ,\unsupported_control_frame_reg[48]_i_1_n_3 ,\unsupported_control_frame_reg[48]_i_1_n_4 ,\unsupported_control_frame_reg[48]_i_1_n_5 ,\unsupported_control_frame_reg[48]_i_1_n_6 ,\unsupported_control_frame_reg[48]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[48]_i_1_n_8 ,\unsupported_control_frame_reg[48]_i_1_n_9 ,\unsupported_control_frame_reg[48]_i_1_n_10 ,\unsupported_control_frame_reg[48]_i_1_n_11 ,\unsupported_control_frame_reg[48]_i_1_n_12 ,\unsupported_control_frame_reg[48]_i_1_n_13 ,\unsupported_control_frame_reg[48]_i_1_n_14 ,\unsupported_control_frame_reg[48]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[55:48]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[49] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[4] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[50] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[51] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[52] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[53] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[54] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[55] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[48]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[56] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[56]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[56]_i_1 
       (.CI(\unsupported_control_frame_reg[48]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_unsupported_control_frame_reg[56]_i_1_CO_UNCONNECTED [7],\unsupported_control_frame_reg[56]_i_1_n_1 ,\unsupported_control_frame_reg[56]_i_1_n_2 ,\unsupported_control_frame_reg[56]_i_1_n_3 ,\unsupported_control_frame_reg[56]_i_1_n_4 ,\unsupported_control_frame_reg[56]_i_1_n_5 ,\unsupported_control_frame_reg[56]_i_1_n_6 ,\unsupported_control_frame_reg[56]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[56]_i_1_n_8 ,\unsupported_control_frame_reg[56]_i_1_n_9 ,\unsupported_control_frame_reg[56]_i_1_n_10 ,\unsupported_control_frame_reg[56]_i_1_n_11 ,\unsupported_control_frame_reg[56]_i_1_n_12 ,\unsupported_control_frame_reg[56]_i_1_n_13 ,\unsupported_control_frame_reg[56]_i_1_n_14 ,\unsupported_control_frame_reg[56]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[63:56]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[57] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[58] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_13 ),
        .Q(unsupported_control_frame_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[59] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_12 ),
        .Q(unsupported_control_frame_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[5] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[60] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_11 ),
        .Q(unsupported_control_frame_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[61] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_10 ),
        .Q(unsupported_control_frame_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[62] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[63] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[56]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[6] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_9 ),
        .Q(unsupported_control_frame_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[7] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[0]_i_1_n_8 ),
        .Q(unsupported_control_frame_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[8] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_15 ),
        .Q(unsupported_control_frame_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \unsupported_control_frame_reg[8]_i_1 
       (.CI(\unsupported_control_frame_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\unsupported_control_frame_reg[8]_i_1_n_0 ,\unsupported_control_frame_reg[8]_i_1_n_1 ,\unsupported_control_frame_reg[8]_i_1_n_2 ,\unsupported_control_frame_reg[8]_i_1_n_3 ,\unsupported_control_frame_reg[8]_i_1_n_4 ,\unsupported_control_frame_reg[8]_i_1_n_5 ,\unsupported_control_frame_reg[8]_i_1_n_6 ,\unsupported_control_frame_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\unsupported_control_frame_reg[8]_i_1_n_8 ,\unsupported_control_frame_reg[8]_i_1_n_9 ,\unsupported_control_frame_reg[8]_i_1_n_10 ,\unsupported_control_frame_reg[8]_i_1_n_11 ,\unsupported_control_frame_reg[8]_i_1_n_12 ,\unsupported_control_frame_reg[8]_i_1_n_13 ,\unsupported_control_frame_reg[8]_i_1_n_14 ,\unsupported_control_frame_reg[8]_i_1_n_15 }),
        .S(unsupported_control_frame_reg[15:8]));
  FDCE #(
    .INIT(1'b0)) 
    \unsupported_control_frame_reg[9] 
       (.C(clk_i),
        .CE(rxStatRegPlus[14]),
        .CLR(rst_i),
        .D(\unsupported_control_frame_reg[8]_i_1_n_14 ),
        .Q(unsupported_control_frame_reg[9]));
endmodule

(* ORIG_REF_NAME = "management_top" *) 
module switch_elements_management_top
   (cfgRxRegData,
    cfgTxRegData,
    mgmt_rd_data,
    CLK,
    in0,
    out,
    \stat_rd_data_reg[63] ,
    \stat_rd_data_reg[63]_0 ,
    clk_i,
    rst_i,
    mgmt_wr_data,
    \recv_config0_reg[0] ,
    mdio_i,
    rxStatRegPlus,
    txStatRegPlus);
  output [52:0]cfgRxRegData;
  output [9:0]cfgTxRegData;
  output [31:0]mgmt_rd_data;
  output CLK;
  output in0;
  input [9:0]out;
  input \stat_rd_data_reg[63] ;
  input \stat_rd_data_reg[63]_0 ;
  input clk_i;
  input rst_i;
  input [31:0]mgmt_wr_data;
  input [0:0]\recv_config0_reg[0] ;
  input mdio_i;
  input [18:0]rxStatRegPlus;
  input [14:0]txStatRegPlus;

  wire CLK;
  wire [52:0]cfgRxRegData;
  wire [9:0]cfgTxRegData;
  wire clk_i;
  wire in0;
  wire [15:0]mdio_data_in;
  wire mdio_i;
  wire mdio_in_valid;
  wire [1:1]mdio_opcode;
  wire mdio_out_valid;
  wire [4:0]mgmt_config;
  wire [31:0]mgmt_rd_data;
  wire [31:0]mgmt_wr_data;
  wire [9:0]out;
  wire [0:0]\recv_config0_reg[0] ;
  wire rst_i;
  wire [18:0]rxStatRegPlus;
  wire \stat_rd_data_reg[63] ;
  wire \stat_rd_data_reg[63]_0 ;
  wire [14:0]txStatRegPlus;

  switch_elements_mdio mdio_inst
       (.Q(mgmt_config),
        .clk_i(clk_i),
        .mdc_reg_0(CLK),
        .\mdio_data_in_reg[15]_0 (mdio_data_in),
        .mdio_i(mdio_i),
        .mdio_in_valid(mdio_in_valid),
        .mdio_opcode(mdio_opcode),
        .mdio_out_valid(mdio_out_valid),
        .rst_i(rst_i));
  switch_elements_manage_registers mgmt_interface
       (.Q(mgmt_config),
        .cfgRxRegData(cfgRxRegData),
        .cfgTxRegData(cfgTxRegData),
        .clk_i(clk_i),
        .in0(in0),
        .mdio_in_valid(mdio_in_valid),
        .mdio_opcode(mdio_opcode),
        .mdio_out_valid(mdio_out_valid),
        .mgmt_rd_data(mgmt_rd_data),
        .\mgmt_rd_data_reg[15]_0 (mdio_data_in),
        .mgmt_wr_data(mgmt_wr_data),
        .out(out),
        .\recv_config0_reg[0]_0 (\recv_config0_reg[0] ),
        .rst_i(rst_i),
        .rxStatRegPlus(rxStatRegPlus),
        .\stat_rd_data_reg[63]_0 (\stat_rd_data_reg[63] ),
        .\stat_rd_data_reg[63]_1 (\stat_rd_data_reg[63]_0 ),
        .txStatRegPlus(txStatRegPlus));
endmodule

(* ORIG_REF_NAME = "manchesterWireless" *) 
module switch_elements_manchesterWireless
   (waitforstart_rdy,
    q_o,
    ready_o,
    in0,
    out,
    clk_i,
    rst_i);
  output waitforstart_rdy;
  output [3:0]q_o;
  output ready_o;
  output [3:0]in0;
  input out;
  input clk_i;
  input rst_i;

  wire clk_i;
  wire double_zero;
  wire [3:0]in0;
  wire inst_decode_n_2;
  wire inst_decode_n_3;
  wire inst_decode_n_4;
  wire inst_decode_n_5;
  wire inst_singleDouble_n_4;
  wire inst_singleDouble_n_5;
  wire inst_singleDouble_n_6;
  wire inst_singleDouble_n_7;
  wire md16_nd;
  wire out;
  wire [3:0]q_o;
  wire q_o11_in;
  wire q_o12_in;
  wire ready_o;
  wire rst_i;
  wire [0:0]state;
  wire waitforstart_rdy;

  switch_elements_decode inst_decode
       (.CO(q_o11_in),
        .D(inst_singleDouble_n_4),
        .\FSM_sequential_state_reg[0]_0 (inst_decode_n_3),
        .\FSM_sequential_state_reg[0]_1 (inst_singleDouble_n_7),
        .\FSM_sequential_state_reg[0]_2 (q_o12_in),
        .\FSM_sequential_state_reg[0]_3 (double_zero),
        .\FSM_sequential_state_reg[1]_0 (inst_decode_n_5),
        .\FSM_sequential_state_reg[2]_0 (inst_decode_n_4),
        .\FSM_sequential_state_reg[2]_1 (inst_singleDouble_n_6),
        .\FSM_sequential_state_reg[2]_2 (inst_singleDouble_n_5),
        .Q(state),
        .clk_i(clk_i),
        .\index_reg[4]_0 (inst_decode_n_2),
        .md16_nd(md16_nd),
        .q_o(q_o),
        .ready_o(ready_o),
        .rst_i(rst_i));
  switch_elements_singleDouble inst_singleDouble
       (.CO(q_o11_in),
        .D(inst_singleDouble_n_4),
        .\FSM_sequential_state_reg[1] (inst_decode_n_2),
        .\FSM_sequential_state_reg[1]_0 (inst_decode_n_5),
        .\FSM_sequential_state_reg[1]_1 (inst_decode_n_4),
        .\FSM_sequential_state_reg[1]_2 (inst_decode_n_3),
        .Q(state),
        .ce_i_d_reg_0(waitforstart_rdy),
        .clk_i(clk_i),
        .\count_zeros_reg[16]_0 (q_o12_in),
        .\count_zeros_reg[16]_1 (double_zero),
        .in0(in0),
        .md16_nd(md16_nd),
        .out(out),
        .rst_i(rst_i),
        .rst_i_0(inst_singleDouble_n_5),
        .rst_i_1(inst_singleDouble_n_6),
        .rst_i_2(inst_singleDouble_n_7));
  switch_elements_waitForStart inst_waitForStart
       (.clk_i(clk_i),
        .out(out),
        .rst_i(rst_i),
        .waitforstart_rdy(waitforstart_rdy));
endmodule

(* ORIG_REF_NAME = "mdio" *) 
module switch_elements_mdio
   (mdc_reg_0,
    mdio_in_valid,
    \mdio_data_in_reg[15]_0 ,
    rst_i,
    clk_i,
    mdio_out_valid,
    mdio_opcode,
    Q,
    mdio_i);
  output mdc_reg_0;
  output mdio_in_valid;
  output [15:0]\mdio_data_in_reg[15]_0 ;
  input rst_i;
  input clk_i;
  input mdio_out_valid;
  input [0:0]mdio_opcode;
  input [4:0]Q;
  input mdio_i;

  wire \FSM_onehot_nextstate_reg[0]_i_1_n_0 ;
  wire \FSM_onehot_nextstate_reg[1]_i_1_n_0 ;
  wire \FSM_onehot_nextstate_reg[2]_i_1_n_0 ;
  wire \FSM_onehot_nextstate_reg_n_0_[0] ;
  wire \FSM_onehot_nextstate_reg_n_0_[1] ;
  wire \FSM_onehot_nextstate_reg_n_0_[2] ;
  wire \FSM_onehot_state_reg_n_0_[0] ;
  wire \FSM_onehot_state_reg_n_0_[1] ;
  wire \FSM_onehot_state_reg_n_0_[2] ;
  wire [4:0]Q;
  wire \clk_cnt[0]_i_1_n_0 ;
  wire \clk_cnt[1]_i_1_n_0 ;
  wire \clk_cnt[2]_i_1_n_0 ;
  wire \clk_cnt[3]_i_1_n_0 ;
  wire \clk_cnt[4]_i_1_n_0 ;
  wire \clk_cnt[4]_i_2_n_0 ;
  wire \clk_cnt[4]_i_3_n_0 ;
  wire [4:0]clk_cnt_reg;
  wire clk_i;
  wire data0;
  wire mdc_i_1_n_0;
  wire mdc_reg_0;
  wire [15:0]\mdio_data_in_reg[15]_0 ;
  wire mdio_i;
  wire mdio_in_valid;
  wire mdio_in_valid_i_2_n_0;
  wire [0:0]mdio_opcode;
  wire mdio_operate_done;
  wire mdio_out_valid;
  wire mdio_t__6;
  wire nextstate;
  wire [6:1]p_0_in;
  wire receiving;
  wire receiving_0;
  wire receiving_i_2_n_0;
  wire receiving_i_5_n_0;
  wire rst_i;
  wire \trans_cnt[0]_i_1_n_0 ;
  wire \trans_cnt[6]_i_2_n_0 ;
  wire [6:0]trans_cnt_reg;
  wire transmitting;
  wire transmitting_1;
  wire transmitting_i_1_n_0;
  wire transmitting_i_3_n_0;
  wire transmitting_i_4_n_0;
  wire transmitting_i_5_n_0;
  wire transmitting_i_6_n_0;

  (* XILINX_LEGACY_PRIM = "LDP" *) 
  LDPE #(
    .INIT(1'b1)) 
    \FSM_onehot_nextstate_reg[0] 
       (.D(\FSM_onehot_nextstate_reg[0]_i_1_n_0 ),
        .G(nextstate),
        .GE(1'b1),
        .PRE(rst_i),
        .Q(\FSM_onehot_nextstate_reg_n_0_[0] ));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hC8)) 
    \FSM_onehot_nextstate_reg[0]_i_1 
       (.I0(\FSM_onehot_state_reg_n_0_[1] ),
        .I1(mdio_operate_done),
        .I2(\FSM_onehot_state_reg_n_0_[2] ),
        .O(\FSM_onehot_nextstate_reg[0]_i_1_n_0 ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_nextstate_reg[1] 
       (.CLR(rst_i),
        .D(\FSM_onehot_nextstate_reg[1]_i_1_n_0 ),
        .G(nextstate),
        .GE(1'b1),
        .Q(\FSM_onehot_nextstate_reg_n_0_[1] ));
  LUT5 #(
    .INIT(32'h20FF2020)) 
    \FSM_onehot_nextstate_reg[1]_i_1 
       (.I0(mdio_out_valid),
        .I1(mdio_opcode),
        .I2(\FSM_onehot_state_reg_n_0_[0] ),
        .I3(mdio_operate_done),
        .I4(\FSM_onehot_state_reg_n_0_[1] ),
        .O(\FSM_onehot_nextstate_reg[1]_i_1_n_0 ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_nextstate_reg[2] 
       (.CLR(rst_i),
        .D(\FSM_onehot_nextstate_reg[2]_i_1_n_0 ),
        .G(nextstate),
        .GE(1'b1),
        .Q(\FSM_onehot_nextstate_reg_n_0_[2] ));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \FSM_onehot_nextstate_reg[2]_i_1 
       (.I0(mdio_out_valid),
        .I1(mdio_opcode),
        .I2(\FSM_onehot_state_reg_n_0_[0] ),
        .I3(mdio_operate_done),
        .I4(\FSM_onehot_state_reg_n_0_[2] ),
        .O(\FSM_onehot_nextstate_reg[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT4 #(
    .INIT(16'hFFEA)) 
    \FSM_onehot_nextstate_reg[2]_i_2 
       (.I0(\FSM_onehot_state_reg_n_0_[2] ),
        .I1(\FSM_onehot_state_reg_n_0_[0] ),
        .I2(mdio_out_valid),
        .I3(\FSM_onehot_state_reg_n_0_[1] ),
        .O(nextstate));
  (* FSM_ENCODED_STATES = "MDIO_WRITE:010,MDIO_READ:100,IDLE:001" *) 
  FDPE #(
    .INIT(1'b1)) 
    \FSM_onehot_state_reg[0] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .D(\FSM_onehot_nextstate_reg_n_0_[0] ),
        .PRE(rst_i),
        .Q(\FSM_onehot_state_reg_n_0_[0] ));
  (* FSM_ENCODED_STATES = "MDIO_WRITE:010,MDIO_READ:100,IDLE:001" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_state_reg[1] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\FSM_onehot_nextstate_reg_n_0_[1] ),
        .Q(\FSM_onehot_state_reg_n_0_[1] ));
  (* FSM_ENCODED_STATES = "MDIO_WRITE:010,MDIO_READ:100,IDLE:001" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_state_reg[2] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\FSM_onehot_nextstate_reg_n_0_[2] ),
        .Q(\FSM_onehot_state_reg_n_0_[2] ));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \clk_cnt[0]_i_1 
       (.I0(clk_cnt_reg[0]),
        .I1(\clk_cnt[4]_i_2_n_0 ),
        .O(\clk_cnt[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \clk_cnt[1]_i_1 
       (.I0(clk_cnt_reg[1]),
        .I1(clk_cnt_reg[0]),
        .I2(\clk_cnt[4]_i_2_n_0 ),
        .O(\clk_cnt[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT4 #(
    .INIT(16'h006A)) 
    \clk_cnt[2]_i_1 
       (.I0(clk_cnt_reg[2]),
        .I1(clk_cnt_reg[1]),
        .I2(clk_cnt_reg[0]),
        .I3(\clk_cnt[4]_i_2_n_0 ),
        .O(\clk_cnt[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'h00006AAA)) 
    \clk_cnt[3]_i_1 
       (.I0(clk_cnt_reg[3]),
        .I1(clk_cnt_reg[2]),
        .I2(clk_cnt_reg[0]),
        .I3(clk_cnt_reg[1]),
        .I4(\clk_cnt[4]_i_2_n_0 ),
        .O(\clk_cnt[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h000000006AAAAAAA)) 
    \clk_cnt[4]_i_1 
       (.I0(clk_cnt_reg[4]),
        .I1(clk_cnt_reg[3]),
        .I2(clk_cnt_reg[1]),
        .I3(clk_cnt_reg[0]),
        .I4(clk_cnt_reg[2]),
        .I5(\clk_cnt[4]_i_2_n_0 ),
        .O(\clk_cnt[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h90000090)) 
    \clk_cnt[4]_i_2 
       (.I0(clk_cnt_reg[3]),
        .I1(Q[3]),
        .I2(\clk_cnt[4]_i_3_n_0 ),
        .I3(Q[4]),
        .I4(clk_cnt_reg[4]),
        .O(\clk_cnt[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \clk_cnt[4]_i_3 
       (.I0(clk_cnt_reg[0]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(clk_cnt_reg[2]),
        .I4(Q[1]),
        .I5(clk_cnt_reg[1]),
        .O(\clk_cnt[4]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \clk_cnt_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\clk_cnt[0]_i_1_n_0 ),
        .Q(clk_cnt_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \clk_cnt_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\clk_cnt[1]_i_1_n_0 ),
        .Q(clk_cnt_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \clk_cnt_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\clk_cnt[2]_i_1_n_0 ),
        .Q(clk_cnt_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \clk_cnt_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\clk_cnt[3]_i_1_n_0 ),
        .Q(clk_cnt_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \clk_cnt_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\clk_cnt[4]_i_1_n_0 ),
        .Q(clk_cnt_reg[4]));
  LUT2 #(
    .INIT(4'h6)) 
    mdc_i_1
       (.I0(\clk_cnt[4]_i_2_n_0 ),
        .I1(mdc_reg_0),
        .O(mdc_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    mdc_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(mdc_i_1_n_0),
        .Q(mdc_reg_0));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[0] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(mdio_i),
        .Q(\mdio_data_in_reg[15]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[10] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [9]),
        .Q(\mdio_data_in_reg[15]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[11] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [10]),
        .Q(\mdio_data_in_reg[15]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[12] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [11]),
        .Q(\mdio_data_in_reg[15]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[13] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [12]),
        .Q(\mdio_data_in_reg[15]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[14] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [13]),
        .Q(\mdio_data_in_reg[15]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[15] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [14]),
        .Q(\mdio_data_in_reg[15]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[1] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [0]),
        .Q(\mdio_data_in_reg[15]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[2] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [1]),
        .Q(\mdio_data_in_reg[15]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[3] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [2]),
        .Q(\mdio_data_in_reg[15]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[4] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [3]),
        .Q(\mdio_data_in_reg[15]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[5] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [4]),
        .Q(\mdio_data_in_reg[15]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[6] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [5]),
        .Q(\mdio_data_in_reg[15]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[7] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [6]),
        .Q(\mdio_data_in_reg[15]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[8] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [7]),
        .Q(\mdio_data_in_reg[15]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \mdio_data_in_reg[9] 
       (.C(mdc_reg_0),
        .CE(receiving),
        .CLR(rst_i),
        .D(\mdio_data_in_reg[15]_0 [8]),
        .Q(\mdio_data_in_reg[15]_0 [9]));
  LUT4 #(
    .INIT(16'h0040)) 
    mdio_in_valid_i_1
       (.I0(trans_cnt_reg[6]),
        .I1(trans_cnt_reg[4]),
        .I2(trans_cnt_reg[5]),
        .I3(mdio_in_valid_i_2_n_0),
        .O(mdio_operate_done));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    mdio_in_valid_i_2
       (.I0(trans_cnt_reg[1]),
        .I1(trans_cnt_reg[0]),
        .I2(trans_cnt_reg[3]),
        .I3(trans_cnt_reg[2]),
        .O(mdio_in_valid_i_2_n_0));
  FDCE #(
    .INIT(1'b0)) 
    mdio_in_valid_reg
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(mdio_operate_done),
        .Q(mdio_in_valid));
  LUT6 #(
    .INIT(64'hAAAAAA2A00000000)) 
    receiving_i_1
       (.I0(\FSM_onehot_state_reg_n_0_[2] ),
        .I1(trans_cnt_reg[5]),
        .I2(trans_cnt_reg[2]),
        .I3(trans_cnt_reg[4]),
        .I4(receiving_i_2_n_0),
        .I5(mdio_t__6),
        .O(receiving_0));
  LUT4 #(
    .INIT(16'hFFF7)) 
    receiving_i_2
       (.I0(trans_cnt_reg[3]),
        .I1(trans_cnt_reg[0]),
        .I2(trans_cnt_reg[1]),
        .I3(trans_cnt_reg[6]),
        .O(receiving_i_2_n_0));
  LUT5 #(
    .INIT(32'hA8AAAAAA)) 
    receiving_i_3
       (.I0(data0),
        .I1(receiving_i_5_n_0),
        .I2(trans_cnt_reg[6]),
        .I3(trans_cnt_reg[0]),
        .I4(trans_cnt_reg[5]),
        .O(mdio_t__6));
  LUT6 #(
    .INIT(64'hFEEEEEEEAAAAAAAA)) 
    receiving_i_4
       (.I0(trans_cnt_reg[6]),
        .I1(trans_cnt_reg[4]),
        .I2(trans_cnt_reg[2]),
        .I3(trans_cnt_reg[3]),
        .I4(trans_cnt_reg[1]),
        .I5(trans_cnt_reg[5]),
        .O(data0));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    receiving_i_5
       (.I0(trans_cnt_reg[3]),
        .I1(trans_cnt_reg[4]),
        .I2(trans_cnt_reg[1]),
        .I3(trans_cnt_reg[2]),
        .O(receiving_i_5_n_0));
  FDCE #(
    .INIT(1'b0)) 
    receiving_reg
       (.C(mdc_reg_0),
        .CE(transmitting_i_1_n_0),
        .CLR(rst_i),
        .D(receiving_0),
        .Q(receiving));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \trans_cnt[0]_i_1 
       (.I0(transmitting),
        .I1(trans_cnt_reg[0]),
        .O(\trans_cnt[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \trans_cnt[1]_i_1 
       (.I0(trans_cnt_reg[1]),
        .I1(trans_cnt_reg[0]),
        .I2(transmitting),
        .O(p_0_in[1]));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT4 #(
    .INIT(16'h6A00)) 
    \trans_cnt[2]_i_1 
       (.I0(trans_cnt_reg[2]),
        .I1(trans_cnt_reg[1]),
        .I2(trans_cnt_reg[0]),
        .I3(transmitting),
        .O(p_0_in[2]));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT5 #(
    .INIT(32'h6AAA0000)) 
    \trans_cnt[3]_i_1 
       (.I0(trans_cnt_reg[3]),
        .I1(trans_cnt_reg[2]),
        .I2(trans_cnt_reg[0]),
        .I3(trans_cnt_reg[1]),
        .I4(transmitting),
        .O(p_0_in[3]));
  LUT6 #(
    .INIT(64'h6AAAAAAA00000000)) 
    \trans_cnt[4]_i_1 
       (.I0(trans_cnt_reg[4]),
        .I1(trans_cnt_reg[3]),
        .I2(trans_cnt_reg[1]),
        .I3(trans_cnt_reg[0]),
        .I4(trans_cnt_reg[2]),
        .I5(transmitting),
        .O(p_0_in[4]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \trans_cnt[5]_i_1 
       (.I0(trans_cnt_reg[5]),
        .I1(\trans_cnt[6]_i_2_n_0 ),
        .I2(transmitting),
        .O(p_0_in[5]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT4 #(
    .INIT(16'h6A00)) 
    \trans_cnt[6]_i_1 
       (.I0(trans_cnt_reg[6]),
        .I1(trans_cnt_reg[5]),
        .I2(\trans_cnt[6]_i_2_n_0 ),
        .I3(transmitting),
        .O(p_0_in[6]));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \trans_cnt[6]_i_2 
       (.I0(trans_cnt_reg[4]),
        .I1(trans_cnt_reg[2]),
        .I2(trans_cnt_reg[0]),
        .I3(trans_cnt_reg[1]),
        .I4(trans_cnt_reg[3]),
        .O(\trans_cnt[6]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[0] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\trans_cnt[0]_i_1_n_0 ),
        .Q(trans_cnt_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[1] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(p_0_in[1]),
        .Q(trans_cnt_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[2] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(p_0_in[2]),
        .Q(trans_cnt_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[3] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(p_0_in[3]),
        .Q(trans_cnt_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[4] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(p_0_in[4]),
        .Q(trans_cnt_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[5] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(p_0_in[5]),
        .Q(trans_cnt_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \trans_cnt_reg[6] 
       (.C(mdc_reg_0),
        .CE(1'b1),
        .CLR(rst_i),
        .D(p_0_in[6]),
        .Q(trans_cnt_reg[6]));
  LUT3 #(
    .INIT(8'hFE)) 
    transmitting_i_1
       (.I0(\FSM_onehot_state_reg_n_0_[1] ),
        .I1(\FSM_onehot_state_reg_n_0_[0] ),
        .I2(\FSM_onehot_state_reg_n_0_[2] ),
        .O(transmitting_i_1_n_0));
  LUT4 #(
    .INIT(16'hFC88)) 
    transmitting_i_2
       (.I0(\FSM_onehot_state_reg_n_0_[1] ),
        .I1(transmitting_i_3_n_0),
        .I2(transmitting_i_4_n_0),
        .I3(\FSM_onehot_state_reg_n_0_[2] ),
        .O(transmitting_1));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'hFFF7)) 
    transmitting_i_3
       (.I0(trans_cnt_reg[5]),
        .I1(trans_cnt_reg[0]),
        .I2(trans_cnt_reg[6]),
        .I3(transmitting_i_5_n_0),
        .O(transmitting_i_3_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    transmitting_i_4
       (.I0(trans_cnt_reg[6]),
        .I1(trans_cnt_reg[4]),
        .I2(trans_cnt_reg[1]),
        .I3(transmitting_i_6_n_0),
        .O(transmitting_i_4_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    transmitting_i_5
       (.I0(trans_cnt_reg[3]),
        .I1(trans_cnt_reg[4]),
        .I2(trans_cnt_reg[1]),
        .I3(trans_cnt_reg[2]),
        .O(transmitting_i_5_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    transmitting_i_6
       (.I0(trans_cnt_reg[2]),
        .I1(trans_cnt_reg[5]),
        .I2(trans_cnt_reg[0]),
        .I3(trans_cnt_reg[3]),
        .O(transmitting_i_6_n_0));
  FDCE #(
    .INIT(1'b0)) 
    transmitting_reg
       (.C(mdc_reg_0),
        .CE(transmitting_i_1_n_0),
        .CLR(rst_i),
        .D(transmitting_1),
        .Q(transmitting));
endmodule

(* ORIG_REF_NAME = "rxCRC" *) 
module switch_elements_rxCRC
   (get_terminator_d1,
    get_terminator_d2,
    get_terminator_d3,
    do_crc_check,
    crc_8_en_reg_0,
    small_error_reg,
    D,
    \bytes_cnt_reg[1]_0 ,
    \bytes_cnt_reg[2]_0 ,
    \CRC_OUT_reg[31] ,
    \CRC_OUT_reg[29] ,
    \CRC_OUT_reg[29]_0 ,
    \CRC_OUT_reg[25] ,
    \rxd64_d3_reg[37] ,
    \CRC_OUT_reg[11] ,
    \CRC_OUT_reg[18] ,
    \rxd64_d3_reg[48] ,
    \CRC_OUT_reg[14] ,
    \CRC_OUT_reg[7] ,
    \CRC_OUT_reg[17] ,
    \CRC_OUT_reg[27] ,
    \rxd64_d3_reg[54] ,
    \CRC_OUT_reg[15] ,
    \CRC_OUT_reg[26] ,
    \CRC_OUT_reg[30] ,
    \CRC_OUT_reg[28] ,
    \CRC_OUT_reg[15]_0 ,
    \CRC_OUT_reg[28]_0 ,
    \CRC_OUT_reg[28]_1 ,
    \CRC_OUT_reg[15]_1 ,
    \CRC_OUT_reg[2] ,
    \CRC_OUT_reg[26]_0 ,
    \rxd64_d3_reg[2] ,
    \rxd64_d3_reg[33] ,
    \CRC_OUT_reg[10] ,
    \CRC_OUT_reg[19] ,
    \CRC_OUT_reg[30]_0 ,
    \CRC_OUT_reg[30]_1 ,
    \CRC_OUT_reg[9] ,
    \CRC_OUT_reg[3] ,
    \CRC_OUT_reg[22] ,
    \CRC_OUT_reg[20] ,
    \CRC_OUT_reg[29]_1 ,
    \CRC_OUT_reg[3]_0 ,
    \CRC_OUT_reg[0] ,
    \CRC_OUT_reg[31]_0 ,
    \CRC_OUT_reg[16] ,
    \rxd64_d3_reg[37]_0 ,
    \CRC_OUT_reg[9]_0 ,
    \CRC_OUT_reg[23] ,
    get_terminator,
    clk_i,
    reset_dcm,
    do_crc_check_reg_0,
    crc_64_en,
    small_error,
    large_error,
    Q,
    wait_crc_check,
    \bytes_cnt_reg[2]_1 ,
    rxd64_d3,
    \CRC_OUT_reg[24] ,
    \CRC_OUT_reg[24]_0 ,
    \CRC_OUT_reg[24]_1 ,
    \CRC_OUT_reg[1] ,
    \CRC_OUT_reg[6] ,
    \CRC_OUT_reg[22]_0 ,
    \CRC_OUT_reg[22]_1 ,
    \CRC_OUT_reg[29]_2 ,
    \CRC_OUT_reg[29]_3 ,
    \CRC_OUT_reg[29]_4 ,
    E,
    \bytes_cnt_reg[1]_1 ,
    SS,
    \CRC_OUT_reg[31]_1 );
  output get_terminator_d1;
  output get_terminator_d2;
  output get_terminator_d3;
  output do_crc_check;
  output crc_8_en_reg_0;
  output small_error_reg;
  output [0:0]D;
  output [1:0]\bytes_cnt_reg[1]_0 ;
  output \bytes_cnt_reg[2]_0 ;
  output [29:0]\CRC_OUT_reg[31] ;
  output \CRC_OUT_reg[29] ;
  output \CRC_OUT_reg[29]_0 ;
  output \CRC_OUT_reg[25] ;
  output \rxd64_d3_reg[37] ;
  output \CRC_OUT_reg[11] ;
  output \CRC_OUT_reg[18] ;
  output \rxd64_d3_reg[48] ;
  output \CRC_OUT_reg[14] ;
  output \CRC_OUT_reg[7] ;
  output \CRC_OUT_reg[17] ;
  output \CRC_OUT_reg[27] ;
  output \rxd64_d3_reg[54] ;
  output \CRC_OUT_reg[15] ;
  output \CRC_OUT_reg[26] ;
  output \CRC_OUT_reg[30] ;
  output \CRC_OUT_reg[28] ;
  output \CRC_OUT_reg[15]_0 ;
  output \CRC_OUT_reg[28]_0 ;
  output \CRC_OUT_reg[28]_1 ;
  output \CRC_OUT_reg[15]_1 ;
  output \CRC_OUT_reg[2] ;
  output \CRC_OUT_reg[26]_0 ;
  output \rxd64_d3_reg[2] ;
  output \rxd64_d3_reg[33] ;
  output \CRC_OUT_reg[10] ;
  output \CRC_OUT_reg[19] ;
  output \CRC_OUT_reg[30]_0 ;
  output \CRC_OUT_reg[30]_1 ;
  output \CRC_OUT_reg[9] ;
  output \CRC_OUT_reg[3] ;
  output \CRC_OUT_reg[22] ;
  output \CRC_OUT_reg[20] ;
  output \CRC_OUT_reg[29]_1 ;
  output \CRC_OUT_reg[3]_0 ;
  output \CRC_OUT_reg[0] ;
  output \CRC_OUT_reg[31]_0 ;
  output \CRC_OUT_reg[16] ;
  output \rxd64_d3_reg[37]_0 ;
  output \CRC_OUT_reg[9]_0 ;
  output \CRC_OUT_reg[23] ;
  input get_terminator;
  input clk_i;
  input reset_dcm;
  input do_crc_check_reg_0;
  input crc_64_en;
  input small_error;
  input large_error;
  input [0:0]Q;
  input wait_crc_check;
  input [0:0]\bytes_cnt_reg[2]_1 ;
  input [63:0]rxd64_d3;
  input \CRC_OUT_reg[24] ;
  input \CRC_OUT_reg[24]_0 ;
  input \CRC_OUT_reg[24]_1 ;
  input \CRC_OUT_reg[1] ;
  input \CRC_OUT_reg[6] ;
  input \CRC_OUT_reg[22]_0 ;
  input \CRC_OUT_reg[22]_1 ;
  input \CRC_OUT_reg[29]_2 ;
  input \CRC_OUT_reg[29]_3 ;
  input \CRC_OUT_reg[29]_4 ;
  input [0:0]E;
  input [1:0]\bytes_cnt_reg[1]_1 ;
  input [0:0]SS;
  input [30:0]\CRC_OUT_reg[31]_1 ;

  wire [7:0]CRC_DATA_TMP;
  wire \CRC_OUT_reg[0] ;
  wire \CRC_OUT_reg[10] ;
  wire \CRC_OUT_reg[11] ;
  wire \CRC_OUT_reg[14] ;
  wire \CRC_OUT_reg[15] ;
  wire \CRC_OUT_reg[15]_0 ;
  wire \CRC_OUT_reg[15]_1 ;
  wire \CRC_OUT_reg[16] ;
  wire \CRC_OUT_reg[17] ;
  wire \CRC_OUT_reg[18] ;
  wire \CRC_OUT_reg[19] ;
  wire \CRC_OUT_reg[1] ;
  wire \CRC_OUT_reg[20] ;
  wire \CRC_OUT_reg[22] ;
  wire \CRC_OUT_reg[22]_0 ;
  wire \CRC_OUT_reg[22]_1 ;
  wire \CRC_OUT_reg[23] ;
  wire \CRC_OUT_reg[24] ;
  wire \CRC_OUT_reg[24]_0 ;
  wire \CRC_OUT_reg[24]_1 ;
  wire \CRC_OUT_reg[25] ;
  wire \CRC_OUT_reg[26] ;
  wire \CRC_OUT_reg[26]_0 ;
  wire \CRC_OUT_reg[27] ;
  wire \CRC_OUT_reg[28] ;
  wire \CRC_OUT_reg[28]_0 ;
  wire \CRC_OUT_reg[28]_1 ;
  wire \CRC_OUT_reg[29] ;
  wire \CRC_OUT_reg[29]_0 ;
  wire \CRC_OUT_reg[29]_1 ;
  wire \CRC_OUT_reg[29]_2 ;
  wire \CRC_OUT_reg[29]_3 ;
  wire \CRC_OUT_reg[29]_4 ;
  wire \CRC_OUT_reg[2] ;
  wire \CRC_OUT_reg[30] ;
  wire \CRC_OUT_reg[30]_0 ;
  wire \CRC_OUT_reg[30]_1 ;
  wire [29:0]\CRC_OUT_reg[31] ;
  wire \CRC_OUT_reg[31]_0 ;
  wire [30:0]\CRC_OUT_reg[31]_1 ;
  wire \CRC_OUT_reg[3] ;
  wire \CRC_OUT_reg[3]_0 ;
  wire \CRC_OUT_reg[6] ;
  wire \CRC_OUT_reg[7] ;
  wire \CRC_OUT_reg[9] ;
  wire \CRC_OUT_reg[9]_0 ;
  wire [0:0]D;
  wire [0:0]E;
  wire [0:0]Q;
  wire [0:0]SS;
  wire [2:2]bytes_cnt;
  wire \bytes_cnt[2]_i_2_n_0 ;
  wire [1:0]\bytes_cnt_reg[1]_0 ;
  wire [1:0]\bytes_cnt_reg[1]_1 ;
  wire \bytes_cnt_reg[2]_0 ;
  wire [0:0]\bytes_cnt_reg[2]_1 ;
  wire clk_i;
  wire crc_64_en;
  wire crc_64_en_reg_n_0;
  wire crc_8_en_i_1_n_0;
  wire crc_8_en_reg_0;
  wire [29:9]crc_from_64;
  wire do_crc_check;
  wire do_crc_check_reg_0;
  wire get_terminator;
  wire get_terminator_d1;
  wire get_terminator_d2;
  wire get_terminator_d3;
  wire large_error;
  wire reset_dcm;
  wire [63:0]rxd64_d3;
  wire \rxd64_d3_reg[2] ;
  wire \rxd64_d3_reg[33] ;
  wire \rxd64_d3_reg[37] ;
  wire \rxd64_d3_reg[37]_0 ;
  wire \rxd64_d3_reg[48] ;
  wire \rxd64_d3_reg[54] ;
  wire small_error;
  wire small_error_reg;
  wire [63:0]terminator_data;
  wire \terminator_data[0]_i_1_n_0 ;
  wire \terminator_data[10]_i_1_n_0 ;
  wire \terminator_data[11]_i_1_n_0 ;
  wire \terminator_data[12]_i_1_n_0 ;
  wire \terminator_data[13]_i_1_n_0 ;
  wire \terminator_data[14]_i_1_n_0 ;
  wire \terminator_data[15]_i_1_n_0 ;
  wire \terminator_data[16]_i_1_n_0 ;
  wire \terminator_data[17]_i_1_n_0 ;
  wire \terminator_data[18]_i_1_n_0 ;
  wire \terminator_data[19]_i_1_n_0 ;
  wire \terminator_data[1]_i_1_n_0 ;
  wire \terminator_data[20]_i_1_n_0 ;
  wire \terminator_data[21]_i_1_n_0 ;
  wire \terminator_data[22]_i_1_n_0 ;
  wire \terminator_data[23]_i_1_n_0 ;
  wire \terminator_data[24]_i_1_n_0 ;
  wire \terminator_data[25]_i_1_n_0 ;
  wire \terminator_data[26]_i_1_n_0 ;
  wire \terminator_data[27]_i_1_n_0 ;
  wire \terminator_data[28]_i_1_n_0 ;
  wire \terminator_data[29]_i_1_n_0 ;
  wire \terminator_data[2]_i_1_n_0 ;
  wire \terminator_data[30]_i_1_n_0 ;
  wire \terminator_data[31]_i_1_n_0 ;
  wire \terminator_data[32]_i_1_n_0 ;
  wire \terminator_data[33]_i_1_n_0 ;
  wire \terminator_data[34]_i_1_n_0 ;
  wire \terminator_data[35]_i_1_n_0 ;
  wire \terminator_data[36]_i_1_n_0 ;
  wire \terminator_data[37]_i_1_n_0 ;
  wire \terminator_data[38]_i_1_n_0 ;
  wire \terminator_data[39]_i_1_n_0 ;
  wire \terminator_data[3]_i_1_n_0 ;
  wire \terminator_data[40]_i_1_n_0 ;
  wire \terminator_data[41]_i_1_n_0 ;
  wire \terminator_data[42]_i_1_n_0 ;
  wire \terminator_data[43]_i_1_n_0 ;
  wire \terminator_data[44]_i_1_n_0 ;
  wire \terminator_data[45]_i_1_n_0 ;
  wire \terminator_data[46]_i_1_n_0 ;
  wire \terminator_data[47]_i_1_n_0 ;
  wire \terminator_data[48]_i_1_n_0 ;
  wire \terminator_data[49]_i_1_n_0 ;
  wire \terminator_data[4]_i_1_n_0 ;
  wire \terminator_data[50]_i_1_n_0 ;
  wire \terminator_data[51]_i_1_n_0 ;
  wire \terminator_data[52]_i_1_n_0 ;
  wire \terminator_data[53]_i_1_n_0 ;
  wire \terminator_data[54]_i_1_n_0 ;
  wire \terminator_data[55]_i_1_n_0 ;
  wire \terminator_data[56]_i_1_n_0 ;
  wire \terminator_data[57]_i_1_n_0 ;
  wire \terminator_data[58]_i_1_n_0 ;
  wire \terminator_data[59]_i_1_n_0 ;
  wire \terminator_data[5]_i_1_n_0 ;
  wire \terminator_data[60]_i_1_n_0 ;
  wire \terminator_data[61]_i_1_n_0 ;
  wire \terminator_data[62]_i_1_n_0 ;
  wire \terminator_data[63]_i_1_n_0 ;
  wire \terminator_data[6]_i_1_n_0 ;
  wire \terminator_data[7]_i_1_n_0 ;
  wire \terminator_data[8]_i_1_n_0 ;
  wire \terminator_data[9]_i_1_n_0 ;
  wire wait_crc_check;

  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[56]),
        .Q(CRC_DATA_TMP[0]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[57]),
        .Q(CRC_DATA_TMP[1]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[58]),
        .Q(CRC_DATA_TMP[2]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[59]),
        .Q(CRC_DATA_TMP[3]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[60]),
        .Q(CRC_DATA_TMP[4]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[61]),
        .Q(CRC_DATA_TMP[5]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[62]),
        .Q(CRC_DATA_TMP[6]));
  FDCE #(
    .INIT(1'b0)) 
    \CRC_DATA_TMP_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(terminator_data[63]),
        .Q(CRC_DATA_TMP[7]));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT5 #(
    .INIT(32'hB8B8B88B)) 
    \bytes_cnt[2]_i_2 
       (.I0(\bytes_cnt_reg[2]_1 ),
        .I1(get_terminator),
        .I2(bytes_cnt),
        .I3(\bytes_cnt_reg[1]_0 [0]),
        .I4(\bytes_cnt_reg[1]_0 [1]),
        .O(\bytes_cnt[2]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \bytes_cnt_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(\bytes_cnt_reg[1]_1 [0]),
        .Q(\bytes_cnt_reg[1]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \bytes_cnt_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(\bytes_cnt_reg[1]_1 [1]),
        .Q(\bytes_cnt_reg[1]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \bytes_cnt_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(\bytes_cnt[2]_i_2_n_0 ),
        .Q(bytes_cnt));
  switch_elements_CRC32_D64_3 crc64
       (.\CRC_OUT_reg[0]_0 (\CRC_OUT_reg[0] ),
        .\CRC_OUT_reg[10]_0 (\CRC_OUT_reg[10] ),
        .\CRC_OUT_reg[11]_0 (\CRC_OUT_reg[11] ),
        .\CRC_OUT_reg[14]_0 (\CRC_OUT_reg[14] ),
        .\CRC_OUT_reg[15]_0 (\CRC_OUT_reg[15] ),
        .\CRC_OUT_reg[15]_1 (\CRC_OUT_reg[15]_0 ),
        .\CRC_OUT_reg[15]_2 (\CRC_OUT_reg[15]_1 ),
        .\CRC_OUT_reg[16]_0 (\CRC_OUT_reg[16] ),
        .\CRC_OUT_reg[17]_0 (\CRC_OUT_reg[17] ),
        .\CRC_OUT_reg[18]_0 (\CRC_OUT_reg[18] ),
        .\CRC_OUT_reg[19]_0 (\CRC_OUT_reg[19] ),
        .\CRC_OUT_reg[1]_0 (\CRC_OUT_reg[1] ),
        .\CRC_OUT_reg[20]_0 (\CRC_OUT_reg[20] ),
        .\CRC_OUT_reg[22]_0 (\CRC_OUT_reg[22] ),
        .\CRC_OUT_reg[22]_1 (\CRC_OUT_reg[22]_0 ),
        .\CRC_OUT_reg[22]_2 (\CRC_OUT_reg[22]_1 ),
        .\CRC_OUT_reg[23]_0 (\CRC_OUT_reg[23] ),
        .\CRC_OUT_reg[24]_0 (\CRC_OUT_reg[24] ),
        .\CRC_OUT_reg[24]_1 (\CRC_OUT_reg[24]_0 ),
        .\CRC_OUT_reg[24]_2 (\CRC_OUT_reg[24]_1 ),
        .\CRC_OUT_reg[25]_0 (\CRC_OUT_reg[25] ),
        .\CRC_OUT_reg[26]_0 (\CRC_OUT_reg[26] ),
        .\CRC_OUT_reg[26]_1 (\CRC_OUT_reg[26]_0 ),
        .\CRC_OUT_reg[27]_0 (\CRC_OUT_reg[27] ),
        .\CRC_OUT_reg[28]_0 (\CRC_OUT_reg[28] ),
        .\CRC_OUT_reg[28]_1 (\CRC_OUT_reg[28]_0 ),
        .\CRC_OUT_reg[28]_2 (\CRC_OUT_reg[28]_1 ),
        .\CRC_OUT_reg[29]_0 (\CRC_OUT_reg[29] ),
        .\CRC_OUT_reg[29]_1 (\CRC_OUT_reg[29]_0 ),
        .\CRC_OUT_reg[29]_2 (\CRC_OUT_reg[29]_1 ),
        .\CRC_OUT_reg[29]_3 (\CRC_OUT_reg[29]_2 ),
        .\CRC_OUT_reg[29]_4 (\CRC_OUT_reg[29]_3 ),
        .\CRC_OUT_reg[29]_5 (\CRC_OUT_reg[29]_4 ),
        .\CRC_OUT_reg[2]_0 (\CRC_OUT_reg[2] ),
        .\CRC_OUT_reg[30]_0 (\CRC_OUT_reg[30] ),
        .\CRC_OUT_reg[30]_1 (\CRC_OUT_reg[30]_0 ),
        .\CRC_OUT_reg[30]_2 (\CRC_OUT_reg[30]_1 ),
        .\CRC_OUT_reg[31]_0 (\CRC_OUT_reg[31]_0 ),
        .\CRC_OUT_reg[31]_1 (\CRC_OUT_reg[31]_1 ),
        .\CRC_OUT_reg[3]_0 (\CRC_OUT_reg[3] ),
        .\CRC_OUT_reg[3]_1 (\CRC_OUT_reg[3]_0 ),
        .\CRC_OUT_reg[6]_0 (\CRC_OUT_reg[6] ),
        .\CRC_OUT_reg[7]_0 (\CRC_OUT_reg[7] ),
        .\CRC_OUT_reg[9]_0 (\CRC_OUT_reg[9] ),
        .\CRC_OUT_reg[9]_1 (\CRC_OUT_reg[9]_0 ),
        .E(crc_64_en_reg_n_0),
        .Q({\CRC_OUT_reg[31] [29:28],crc_from_64[29],\CRC_OUT_reg[31] [27:9],crc_from_64[9],\CRC_OUT_reg[31] [8:0]}),
        .SS(SS),
        .clk_i(clk_i),
        .rxd64_d3({rxd64_d3[54],rxd64_d3[49:48],rxd64_d3[39:35],rxd64_d3[33],rxd64_d3[31],rxd64_d3[29:27],rxd64_d3[24],rxd64_d3[22:0]}),
        .\rxd64_d3_reg[2] (\rxd64_d3_reg[2] ),
        .\rxd64_d3_reg[33] (\rxd64_d3_reg[33] ),
        .\rxd64_d3_reg[37] (\rxd64_d3_reg[37] ),
        .\rxd64_d3_reg[37]_0 (\rxd64_d3_reg[37]_0 ),
        .\rxd64_d3_reg[48] (\rxd64_d3_reg[48] ),
        .\rxd64_d3_reg[54] (\rxd64_d3_reg[54] ));
  switch_elements_CRC32_D8_4 crc8
       (.\CRC_OUT_reg[19]_0 (crc_8_en_reg_0),
        .\CRC_OUT_reg[30]_0 (CRC_DATA_TMP),
        .\CRC_OUT_reg[31]_0 ({\CRC_OUT_reg[31] [29:28],crc_from_64[29],\CRC_OUT_reg[31] [27:9],crc_from_64[9],\CRC_OUT_reg[31] [8:0]}),
        .D(D),
        .Q(Q),
        .clk_i(clk_i),
        .do_crc_check(do_crc_check),
        .large_error(large_error),
        .reset_dcm(reset_dcm),
        .small_error(small_error),
        .small_error_reg(small_error_reg),
        .wait_crc_check(wait_crc_check));
  FDCE #(
    .INIT(1'b0)) 
    crc_64_en_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(crc_64_en),
        .Q(crc_64_en_reg_n_0));
  LUT5 #(
    .INIT(32'hFFEFAAAA)) 
    crc_8_en_i_1
       (.I0(get_terminator_d3),
        .I1(\bytes_cnt_reg[1]_0 [1]),
        .I2(\bytes_cnt_reg[1]_0 [0]),
        .I3(bytes_cnt),
        .I4(crc_8_en_reg_0),
        .O(crc_8_en_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    crc_8_en_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(crc_8_en_i_1_n_0),
        .Q(crc_8_en_reg_0));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'h04)) 
    do_crc_check_i_2
       (.I0(bytes_cnt),
        .I1(\bytes_cnt_reg[1]_0 [0]),
        .I2(\bytes_cnt_reg[1]_0 [1]),
        .O(\bytes_cnt_reg[2]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    do_crc_check_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(do_crc_check_reg_0),
        .Q(do_crc_check));
  FDCE #(
    .INIT(1'b0)) 
    get_terminator_d1_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(get_terminator),
        .Q(get_terminator_d1));
  FDCE #(
    .INIT(1'b0)) 
    get_terminator_d2_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(get_terminator_d1),
        .Q(get_terminator_d2));
  FDCE #(
    .INIT(1'b0)) 
    get_terminator_d3_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(get_terminator_d2),
        .Q(get_terminator_d3));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[0]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[63]),
        .O(\terminator_data[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[10]_i_1 
       (.I0(rxd64_d3[53]),
        .I1(get_terminator_d2),
        .I2(terminator_data[2]),
        .O(\terminator_data[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[11]_i_1 
       (.I0(rxd64_d3[52]),
        .I1(get_terminator_d2),
        .I2(terminator_data[3]),
        .O(\terminator_data[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[12]_i_1 
       (.I0(rxd64_d3[51]),
        .I1(get_terminator_d2),
        .I2(terminator_data[4]),
        .O(\terminator_data[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[13]_i_1 
       (.I0(rxd64_d3[50]),
        .I1(get_terminator_d2),
        .I2(terminator_data[5]),
        .O(\terminator_data[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[14]_i_1 
       (.I0(rxd64_d3[49]),
        .I1(get_terminator_d2),
        .I2(terminator_data[6]),
        .O(\terminator_data[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[15]_i_1 
       (.I0(rxd64_d3[48]),
        .I1(get_terminator_d2),
        .I2(terminator_data[7]),
        .O(\terminator_data[15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[16]_i_1 
       (.I0(rxd64_d3[47]),
        .I1(get_terminator_d2),
        .I2(terminator_data[8]),
        .O(\terminator_data[16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[17]_i_1 
       (.I0(rxd64_d3[46]),
        .I1(get_terminator_d2),
        .I2(terminator_data[9]),
        .O(\terminator_data[17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[18]_i_1 
       (.I0(rxd64_d3[45]),
        .I1(get_terminator_d2),
        .I2(terminator_data[10]),
        .O(\terminator_data[18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[19]_i_1 
       (.I0(rxd64_d3[44]),
        .I1(get_terminator_d2),
        .I2(terminator_data[11]),
        .O(\terminator_data[19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[1]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[62]),
        .O(\terminator_data[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[20]_i_1 
       (.I0(rxd64_d3[43]),
        .I1(get_terminator_d2),
        .I2(terminator_data[12]),
        .O(\terminator_data[20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[21]_i_1 
       (.I0(rxd64_d3[42]),
        .I1(get_terminator_d2),
        .I2(terminator_data[13]),
        .O(\terminator_data[21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[22]_i_1 
       (.I0(rxd64_d3[41]),
        .I1(get_terminator_d2),
        .I2(terminator_data[14]),
        .O(\terminator_data[22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[23]_i_1 
       (.I0(rxd64_d3[40]),
        .I1(get_terminator_d2),
        .I2(terminator_data[15]),
        .O(\terminator_data[23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[24]_i_1 
       (.I0(rxd64_d3[39]),
        .I1(get_terminator_d2),
        .I2(terminator_data[16]),
        .O(\terminator_data[24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[25]_i_1 
       (.I0(rxd64_d3[38]),
        .I1(get_terminator_d2),
        .I2(terminator_data[17]),
        .O(\terminator_data[25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[26]_i_1 
       (.I0(rxd64_d3[37]),
        .I1(get_terminator_d2),
        .I2(terminator_data[18]),
        .O(\terminator_data[26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[27]_i_1 
       (.I0(rxd64_d3[36]),
        .I1(get_terminator_d2),
        .I2(terminator_data[19]),
        .O(\terminator_data[27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[28]_i_1 
       (.I0(rxd64_d3[35]),
        .I1(get_terminator_d2),
        .I2(terminator_data[20]),
        .O(\terminator_data[28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[29]_i_1 
       (.I0(rxd64_d3[34]),
        .I1(get_terminator_d2),
        .I2(terminator_data[21]),
        .O(\terminator_data[29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[2]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[61]),
        .O(\terminator_data[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[30]_i_1 
       (.I0(rxd64_d3[33]),
        .I1(get_terminator_d2),
        .I2(terminator_data[22]),
        .O(\terminator_data[30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[31]_i_1 
       (.I0(rxd64_d3[32]),
        .I1(get_terminator_d2),
        .I2(terminator_data[23]),
        .O(\terminator_data[31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[32]_i_1 
       (.I0(rxd64_d3[31]),
        .I1(get_terminator_d2),
        .I2(terminator_data[24]),
        .O(\terminator_data[32]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[33]_i_1 
       (.I0(rxd64_d3[30]),
        .I1(get_terminator_d2),
        .I2(terminator_data[25]),
        .O(\terminator_data[33]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[34]_i_1 
       (.I0(rxd64_d3[29]),
        .I1(get_terminator_d2),
        .I2(terminator_data[26]),
        .O(\terminator_data[34]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[35]_i_1 
       (.I0(rxd64_d3[28]),
        .I1(get_terminator_d2),
        .I2(terminator_data[27]),
        .O(\terminator_data[35]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[36]_i_1 
       (.I0(rxd64_d3[27]),
        .I1(get_terminator_d2),
        .I2(terminator_data[28]),
        .O(\terminator_data[36]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[37]_i_1 
       (.I0(rxd64_d3[26]),
        .I1(get_terminator_d2),
        .I2(terminator_data[29]),
        .O(\terminator_data[37]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[38]_i_1 
       (.I0(rxd64_d3[25]),
        .I1(get_terminator_d2),
        .I2(terminator_data[30]),
        .O(\terminator_data[38]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[39]_i_1 
       (.I0(rxd64_d3[24]),
        .I1(get_terminator_d2),
        .I2(terminator_data[31]),
        .O(\terminator_data[39]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[3]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[60]),
        .O(\terminator_data[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[40]_i_1 
       (.I0(rxd64_d3[23]),
        .I1(get_terminator_d2),
        .I2(terminator_data[32]),
        .O(\terminator_data[40]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[41]_i_1 
       (.I0(rxd64_d3[22]),
        .I1(get_terminator_d2),
        .I2(terminator_data[33]),
        .O(\terminator_data[41]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[42]_i_1 
       (.I0(rxd64_d3[21]),
        .I1(get_terminator_d2),
        .I2(terminator_data[34]),
        .O(\terminator_data[42]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[43]_i_1 
       (.I0(rxd64_d3[20]),
        .I1(get_terminator_d2),
        .I2(terminator_data[35]),
        .O(\terminator_data[43]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[44]_i_1 
       (.I0(rxd64_d3[19]),
        .I1(get_terminator_d2),
        .I2(terminator_data[36]),
        .O(\terminator_data[44]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[45]_i_1 
       (.I0(rxd64_d3[18]),
        .I1(get_terminator_d2),
        .I2(terminator_data[37]),
        .O(\terminator_data[45]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[46]_i_1 
       (.I0(rxd64_d3[17]),
        .I1(get_terminator_d2),
        .I2(terminator_data[38]),
        .O(\terminator_data[46]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[47]_i_1 
       (.I0(rxd64_d3[16]),
        .I1(get_terminator_d2),
        .I2(terminator_data[39]),
        .O(\terminator_data[47]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[48]_i_1 
       (.I0(rxd64_d3[15]),
        .I1(get_terminator_d2),
        .I2(terminator_data[40]),
        .O(\terminator_data[48]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[49]_i_1 
       (.I0(rxd64_d3[14]),
        .I1(get_terminator_d2),
        .I2(terminator_data[41]),
        .O(\terminator_data[49]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[4]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[59]),
        .O(\terminator_data[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[50]_i_1 
       (.I0(rxd64_d3[13]),
        .I1(get_terminator_d2),
        .I2(terminator_data[42]),
        .O(\terminator_data[50]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[51]_i_1 
       (.I0(rxd64_d3[12]),
        .I1(get_terminator_d2),
        .I2(terminator_data[43]),
        .O(\terminator_data[51]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[52]_i_1 
       (.I0(rxd64_d3[11]),
        .I1(get_terminator_d2),
        .I2(terminator_data[44]),
        .O(\terminator_data[52]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[53]_i_1 
       (.I0(rxd64_d3[10]),
        .I1(get_terminator_d2),
        .I2(terminator_data[45]),
        .O(\terminator_data[53]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[54]_i_1 
       (.I0(rxd64_d3[9]),
        .I1(get_terminator_d2),
        .I2(terminator_data[46]),
        .O(\terminator_data[54]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[55]_i_1 
       (.I0(rxd64_d3[8]),
        .I1(get_terminator_d2),
        .I2(terminator_data[47]),
        .O(\terminator_data[55]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[56]_i_1 
       (.I0(rxd64_d3[7]),
        .I1(get_terminator_d2),
        .I2(terminator_data[48]),
        .O(\terminator_data[56]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[57]_i_1 
       (.I0(rxd64_d3[6]),
        .I1(get_terminator_d2),
        .I2(terminator_data[49]),
        .O(\terminator_data[57]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[58]_i_1 
       (.I0(rxd64_d3[5]),
        .I1(get_terminator_d2),
        .I2(terminator_data[50]),
        .O(\terminator_data[58]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[59]_i_1 
       (.I0(rxd64_d3[4]),
        .I1(get_terminator_d2),
        .I2(terminator_data[51]),
        .O(\terminator_data[59]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[5]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[58]),
        .O(\terminator_data[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[60]_i_1 
       (.I0(rxd64_d3[3]),
        .I1(get_terminator_d2),
        .I2(terminator_data[52]),
        .O(\terminator_data[60]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[61]_i_1 
       (.I0(rxd64_d3[2]),
        .I1(get_terminator_d2),
        .I2(terminator_data[53]),
        .O(\terminator_data[61]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[62]_i_1 
       (.I0(rxd64_d3[1]),
        .I1(get_terminator_d2),
        .I2(terminator_data[54]),
        .O(\terminator_data[62]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[63]_i_1 
       (.I0(rxd64_d3[0]),
        .I1(get_terminator_d2),
        .I2(terminator_data[55]),
        .O(\terminator_data[63]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[6]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[57]),
        .O(\terminator_data[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \terminator_data[7]_i_1 
       (.I0(get_terminator_d2),
        .I1(rxd64_d3[56]),
        .O(\terminator_data[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[8]_i_1 
       (.I0(rxd64_d3[55]),
        .I1(get_terminator_d2),
        .I2(terminator_data[0]),
        .O(\terminator_data[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \terminator_data[9]_i_1 
       (.I0(rxd64_d3[54]),
        .I1(get_terminator_d2),
        .I2(terminator_data[1]),
        .O(\terminator_data[9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[0]_i_1_n_0 ),
        .Q(terminator_data[0]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[10]_i_1_n_0 ),
        .Q(terminator_data[10]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[11]_i_1_n_0 ),
        .Q(terminator_data[11]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[12]_i_1_n_0 ),
        .Q(terminator_data[12]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[13]_i_1_n_0 ),
        .Q(terminator_data[13]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[14]_i_1_n_0 ),
        .Q(terminator_data[14]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[15]_i_1_n_0 ),
        .Q(terminator_data[15]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[16]_i_1_n_0 ),
        .Q(terminator_data[16]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[17]_i_1_n_0 ),
        .Q(terminator_data[17]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[18]_i_1_n_0 ),
        .Q(terminator_data[18]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[19]_i_1_n_0 ),
        .Q(terminator_data[19]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[1]_i_1_n_0 ),
        .Q(terminator_data[1]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[20]_i_1_n_0 ),
        .Q(terminator_data[20]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[21]_i_1_n_0 ),
        .Q(terminator_data[21]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[22]_i_1_n_0 ),
        .Q(terminator_data[22]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[23]_i_1_n_0 ),
        .Q(terminator_data[23]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[24]_i_1_n_0 ),
        .Q(terminator_data[24]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[25]_i_1_n_0 ),
        .Q(terminator_data[25]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[26]_i_1_n_0 ),
        .Q(terminator_data[26]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[27]_i_1_n_0 ),
        .Q(terminator_data[27]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[28]_i_1_n_0 ),
        .Q(terminator_data[28]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[29]_i_1_n_0 ),
        .Q(terminator_data[29]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[2]_i_1_n_0 ),
        .Q(terminator_data[2]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[30]_i_1_n_0 ),
        .Q(terminator_data[30]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[31]_i_1_n_0 ),
        .Q(terminator_data[31]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[32]_i_1_n_0 ),
        .Q(terminator_data[32]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[33]_i_1_n_0 ),
        .Q(terminator_data[33]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[34]_i_1_n_0 ),
        .Q(terminator_data[34]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[35]_i_1_n_0 ),
        .Q(terminator_data[35]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[36]_i_1_n_0 ),
        .Q(terminator_data[36]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[37]_i_1_n_0 ),
        .Q(terminator_data[37]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[38]_i_1_n_0 ),
        .Q(terminator_data[38]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[39]_i_1_n_0 ),
        .Q(terminator_data[39]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[3]_i_1_n_0 ),
        .Q(terminator_data[3]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[40]_i_1_n_0 ),
        .Q(terminator_data[40]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[41]_i_1_n_0 ),
        .Q(terminator_data[41]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[42]_i_1_n_0 ),
        .Q(terminator_data[42]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[43]_i_1_n_0 ),
        .Q(terminator_data[43]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[44]_i_1_n_0 ),
        .Q(terminator_data[44]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[45]_i_1_n_0 ),
        .Q(terminator_data[45]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[46]_i_1_n_0 ),
        .Q(terminator_data[46]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[47]_i_1_n_0 ),
        .Q(terminator_data[47]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[48]_i_1_n_0 ),
        .Q(terminator_data[48]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[49]_i_1_n_0 ),
        .Q(terminator_data[49]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[4]_i_1_n_0 ),
        .Q(terminator_data[4]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[50]_i_1_n_0 ),
        .Q(terminator_data[50]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[51]_i_1_n_0 ),
        .Q(terminator_data[51]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[52]_i_1_n_0 ),
        .Q(terminator_data[52]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[53]_i_1_n_0 ),
        .Q(terminator_data[53]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[54]_i_1_n_0 ),
        .Q(terminator_data[54]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[55]_i_1_n_0 ),
        .Q(terminator_data[55]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[56]_i_1_n_0 ),
        .Q(terminator_data[56]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[57]_i_1_n_0 ),
        .Q(terminator_data[57]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[58]_i_1_n_0 ),
        .Q(terminator_data[58]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[59]_i_1_n_0 ),
        .Q(terminator_data[59]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[5]_i_1_n_0 ),
        .Q(terminator_data[5]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[60]_i_1_n_0 ),
        .Q(terminator_data[60]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[61]_i_1_n_0 ),
        .Q(terminator_data[61]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[62]_i_1_n_0 ),
        .Q(terminator_data[62]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[63]_i_1_n_0 ),
        .Q(terminator_data[63]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[6]_i_1_n_0 ),
        .Q(terminator_data[6]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[7]_i_1_n_0 ),
        .Q(terminator_data[7]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[8]_i_1_n_0 ),
        .Q(terminator_data[8]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_data_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\terminator_data[9]_i_1_n_0 ),
        .Q(terminator_data[9]));
endmodule

(* ORIG_REF_NAME = "rxDAchecker" *) 
module switch_elements_rxDAchecker
   (broad_valid,
    multi_valid,
    broad_valid_reg_0,
    clk_i,
    reset_dcm,
    multi_valid_reg_0);
  output broad_valid;
  output multi_valid;
  input broad_valid_reg_0;
  input clk_i;
  input reset_dcm;
  input multi_valid_reg_0;

  wire broad_valid;
  wire broad_valid_reg_0;
  wire clk_i;
  wire multi_valid;
  wire multi_valid_reg_0;
  wire reset_dcm;

  FDCE #(
    .INIT(1'b0)) 
    broad_valid_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(broad_valid_reg_0),
        .Q(broad_valid));
  FDCE #(
    .INIT(1'b0)) 
    multi_valid_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(multi_valid_reg_0),
        .Q(multi_valid));
endmodule

(* ORIG_REF_NAME = "rxDataPath" *) 
module switch_elements_rxDataPath
   (get_error_code,
    get_sfd,
    get_terminator,
    tagged_frame,
    check_reset,
    in0,
    rxd64_d3,
    \FSM_sequential_fifo_state_reg[0]_0 ,
    bad_frame_get_reg,
    good_frame_get_reg,
    get_terminator_reg_0,
    \terminator_location_reg[1]_0 ,
    \terminator_location_reg[2]_0 ,
    get_terminator_d2_reg,
    SS,
    \CRC_OUT_reg[27] ,
    \rxd64_d3_reg[30]_0 ,
    \rxd64_d3_reg[20]_0 ,
    \rxd64_d3_reg[34]_0 ,
    \CRC_OUT_reg[6] ,
    \CRC_OUT_reg[5] ,
    \rxd64_d3_reg[29]_0 ,
    \CRC_OUT_reg[18] ,
    \rxd64_d3_reg[8]_0 ,
    \rxd64_d3_reg[40]_0 ,
    \rxd64_d3_reg[9]_0 ,
    \rx_data_valid_reg[7]_0 ,
    \rx_data_reg[63]_0 ,
    \da_addr_reg[6]_0 ,
    \da_addr_reg[40]_0 ,
    clk_i,
    reset_dcm,
    get_sfd0,
    E,
    Q,
    tagged_frame_reg_0,
    check_reset_reg_0,
    receiving,
    this_cycle,
    get_error_code_reg_0,
    get_terminator_d1,
    bad_frame_get,
    good_frame_get,
    \bytes_cnt_reg[2] ,
    \bytes_cnt_reg[1] ,
    get_terminator_d2,
    wait_crc_check,
    do_crc_check_reg,
    get_terminator_d3,
    rst_i,
    recv_rst,
    \CRC_OUT_reg[11] ,
    \CRC_OUT_reg[1] ,
    \CRC_OUT_reg[10] ,
    \CRC_OUT_reg[13] ,
    \CRC_OUT_reg[24] ,
    \CRC_OUT_reg[24]_0 ,
    \CRC_OUT_reg[6]_0 ,
    \CRC_OUT_reg[6]_1 ,
    \CRC_OUT_reg[28] ,
    \CRC_OUT_reg[28]_0 ,
    \CRC_OUT_reg[26] ,
    \CRC_OUT_reg[9] ,
    \CRC_OUT_reg[9]_0 ,
    \CRC_OUT_reg[22] ,
    \CRC_OUT_reg[30] ,
    \CRC_OUT_reg[14] ,
    \CRC_OUT_reg[31] ,
    \CRC_OUT_reg[9]_1 ,
    \CRC_OUT_reg[18]_0 ,
    \CRC_OUT_reg[18]_1 ,
    \CRC_OUT_reg[8] ,
    \CRC_OUT_reg[8]_0 ,
    \CRC_OUT_reg[16] ,
    \CRC_OUT_reg[5]_0 ,
    \CRC_OUT_reg[5]_1 ,
    \CRC_OUT_reg[1]_0 ,
    \CRC_OUT_reg[12] ,
    \CRC_OUT_reg[20] ,
    \CRC_OUT_reg[23] ,
    \CRC_OUT_reg[13]_0 ,
    \CRC_OUT_reg[15] ,
    \CRC_OUT_reg[15]_0 ,
    \CRC_OUT_reg[17] ,
    \CRC_OUT_reg[14]_0 ,
    \CRC_OUT_reg[25] ,
    \CRC_OUT_reg[22]_0 ,
    \CRC_OUT_reg[4] ,
    \CRC_OUT_reg[8]_1 ,
    \CRC_OUT_reg[8]_2 ,
    \CRC_OUT_reg[11]_0 ,
    \CRC_OUT_reg[18]_2 ,
    qvDataOut,
    D,
    \get_e_chk_reg[7]_0 ,
    \terminator_location_reg[2]_1 ,
    inband_fcs);
  output get_error_code;
  output get_sfd;
  output get_terminator;
  output tagged_frame;
  output check_reset;
  output [0:0]in0;
  output [63:0]rxd64_d3;
  output [0:0]\FSM_sequential_fifo_state_reg[0]_0 ;
  output bad_frame_get_reg;
  output good_frame_get_reg;
  output [0:0]get_terminator_reg_0;
  output [1:0]\terminator_location_reg[1]_0 ;
  output [2:0]\terminator_location_reg[2]_0 ;
  output get_terminator_d2_reg;
  output [0:0]SS;
  output [30:0]\CRC_OUT_reg[27] ;
  output \rxd64_d3_reg[30]_0 ;
  output \rxd64_d3_reg[20]_0 ;
  output \rxd64_d3_reg[34]_0 ;
  output \CRC_OUT_reg[6] ;
  output \CRC_OUT_reg[5] ;
  output \rxd64_d3_reg[29]_0 ;
  output \CRC_OUT_reg[18] ;
  output \rxd64_d3_reg[8]_0 ;
  output \rxd64_d3_reg[40]_0 ;
  output \rxd64_d3_reg[9]_0 ;
  output [7:0]\rx_data_valid_reg[7]_0 ;
  output [63:0]\rx_data_reg[63]_0 ;
  output \da_addr_reg[6]_0 ;
  output \da_addr_reg[40]_0 ;
  input clk_i;
  input reset_dcm;
  input get_sfd0;
  input [0:0]E;
  input [1:0]Q;
  input tagged_frame_reg_0;
  input check_reset_reg_0;
  input receiving;
  input this_cycle;
  input get_error_code_reg_0;
  input get_terminator_d1;
  input bad_frame_get;
  input good_frame_get;
  input \bytes_cnt_reg[2] ;
  input [1:0]\bytes_cnt_reg[1] ;
  input get_terminator_d2;
  input wait_crc_check;
  input do_crc_check_reg;
  input get_terminator_d3;
  input rst_i;
  input recv_rst;
  input \CRC_OUT_reg[11] ;
  input [29:0]\CRC_OUT_reg[1] ;
  input \CRC_OUT_reg[10] ;
  input \CRC_OUT_reg[13] ;
  input \CRC_OUT_reg[24] ;
  input \CRC_OUT_reg[24]_0 ;
  input \CRC_OUT_reg[6]_0 ;
  input \CRC_OUT_reg[6]_1 ;
  input \CRC_OUT_reg[28] ;
  input \CRC_OUT_reg[28]_0 ;
  input \CRC_OUT_reg[26] ;
  input \CRC_OUT_reg[9] ;
  input \CRC_OUT_reg[9]_0 ;
  input \CRC_OUT_reg[22] ;
  input \CRC_OUT_reg[30] ;
  input \CRC_OUT_reg[14] ;
  input \CRC_OUT_reg[31] ;
  input \CRC_OUT_reg[9]_1 ;
  input \CRC_OUT_reg[18]_0 ;
  input \CRC_OUT_reg[18]_1 ;
  input \CRC_OUT_reg[8] ;
  input \CRC_OUT_reg[8]_0 ;
  input \CRC_OUT_reg[16] ;
  input \CRC_OUT_reg[5]_0 ;
  input \CRC_OUT_reg[5]_1 ;
  input \CRC_OUT_reg[1]_0 ;
  input \CRC_OUT_reg[12] ;
  input \CRC_OUT_reg[20] ;
  input \CRC_OUT_reg[23] ;
  input \CRC_OUT_reg[13]_0 ;
  input \CRC_OUT_reg[15] ;
  input \CRC_OUT_reg[15]_0 ;
  input \CRC_OUT_reg[17] ;
  input \CRC_OUT_reg[14]_0 ;
  input \CRC_OUT_reg[25] ;
  input \CRC_OUT_reg[22]_0 ;
  input \CRC_OUT_reg[4] ;
  input \CRC_OUT_reg[8]_1 ;
  input \CRC_OUT_reg[8]_2 ;
  input \CRC_OUT_reg[11]_0 ;
  input \CRC_OUT_reg[18]_2 ;
  input [71:0]qvDataOut;
  input [5:0]D;
  input [7:0]\get_e_chk_reg[7]_0 ;
  input [2:0]\terminator_location_reg[2]_1 ;
  input inband_fcs;

  wire \CRC_OUT[0]_i_2_n_0 ;
  wire \CRC_OUT[0]_i_3_n_0 ;
  wire \CRC_OUT[0]_i_4_n_0 ;
  wire \CRC_OUT[10]_i_2_n_0 ;
  wire \CRC_OUT[10]_i_3_n_0 ;
  wire \CRC_OUT[10]_i_5_n_0 ;
  wire \CRC_OUT[11]_i_2_n_0 ;
  wire \CRC_OUT[11]_i_3_n_0 ;
  wire \CRC_OUT[11]_i_4_n_0 ;
  wire \CRC_OUT[11]_i_5_n_0 ;
  wire \CRC_OUT[11]_i_6_n_0 ;
  wire \CRC_OUT[12]_i_2_n_0 ;
  wire \CRC_OUT[12]_i_3_n_0 ;
  wire \CRC_OUT[13]_i_2_n_0 ;
  wire \CRC_OUT[13]_i_3_n_0 ;
  wire \CRC_OUT[13]_i_4_n_0 ;
  wire \CRC_OUT[13]_i_5_n_0 ;
  wire \CRC_OUT[13]_i_6_n_0 ;
  wire \CRC_OUT[14]_i_2_n_0 ;
  wire \CRC_OUT[14]_i_3_n_0 ;
  wire \CRC_OUT[14]_i_4_n_0 ;
  wire \CRC_OUT[14]_i_5_n_0 ;
  wire \CRC_OUT[15]_i_2_n_0 ;
  wire \CRC_OUT[15]_i_3_n_0 ;
  wire \CRC_OUT[15]_i_4_n_0 ;
  wire \CRC_OUT[16]_i_2_n_0 ;
  wire \CRC_OUT[16]_i_3_n_0 ;
  wire \CRC_OUT[16]_i_4_n_0 ;
  wire \CRC_OUT[16]_i_5_n_0 ;
  wire \CRC_OUT[17]_i_2_n_0 ;
  wire \CRC_OUT[17]_i_3_n_0 ;
  wire \CRC_OUT[17]_i_4_n_0 ;
  wire \CRC_OUT[17]_i_6_n_0 ;
  wire \CRC_OUT[18]_i_2_n_0 ;
  wire \CRC_OUT[18]_i_3_n_0 ;
  wire \CRC_OUT[19]_i_2_n_0 ;
  wire \CRC_OUT[19]_i_3_n_0 ;
  wire \CRC_OUT[19]_i_5_n_0 ;
  wire \CRC_OUT[19]_i_6_n_0 ;
  wire \CRC_OUT[1]_i_2_n_0 ;
  wire \CRC_OUT[1]_i_3_n_0 ;
  wire \CRC_OUT[20]_i_2_n_0 ;
  wire \CRC_OUT[20]_i_3_n_0 ;
  wire \CRC_OUT[20]_i_4_n_0 ;
  wire \CRC_OUT[20]_i_5_n_0 ;
  wire \CRC_OUT[21]_i_2_n_0 ;
  wire \CRC_OUT[21]_i_3_n_0 ;
  wire \CRC_OUT[21]_i_4_n_0 ;
  wire \CRC_OUT[22]_i_2_n_0 ;
  wire \CRC_OUT[22]_i_4_n_0 ;
  wire \CRC_OUT[22]_i_5_n_0 ;
  wire \CRC_OUT[22]_i_6_n_0 ;
  wire \CRC_OUT[23]_i_2_n_0 ;
  wire \CRC_OUT[23]_i_4_n_0 ;
  wire \CRC_OUT[23]_i_5_n_0 ;
  wire \CRC_OUT[23]_i_6_n_0 ;
  wire \CRC_OUT[24]_i_2_n_0 ;
  wire \CRC_OUT[24]_i_3_n_0 ;
  wire \CRC_OUT[24]_i_4_n_0 ;
  wire \CRC_OUT[24]_i_6_n_0 ;
  wire \CRC_OUT[24]_i_8_n_0 ;
  wire \CRC_OUT[25]_i_10_n_0 ;
  wire \CRC_OUT[25]_i_2_n_0 ;
  wire \CRC_OUT[25]_i_3_n_0 ;
  wire \CRC_OUT[25]_i_4_n_0 ;
  wire \CRC_OUT[25]_i_6_n_0 ;
  wire \CRC_OUT[25]_i_8_n_0 ;
  wire \CRC_OUT[25]_i_9_n_0 ;
  wire \CRC_OUT[26]_i_2_n_0 ;
  wire \CRC_OUT[26]_i_4_n_0 ;
  wire \CRC_OUT[26]_i_5_n_0 ;
  wire \CRC_OUT[26]_i_6_n_0 ;
  wire \CRC_OUT[26]_i_7_n_0 ;
  wire \CRC_OUT[26]_i_8_n_0 ;
  wire \CRC_OUT[27]_i_2_n_0 ;
  wire \CRC_OUT[27]_i_4_n_0 ;
  wire \CRC_OUT[27]_i_5_n_0 ;
  wire \CRC_OUT[27]_i_6_n_0 ;
  wire \CRC_OUT[27]_i_7_n_0 ;
  wire \CRC_OUT[27]_i_8_n_0 ;
  wire \CRC_OUT[28]_i_10_n_0 ;
  wire \CRC_OUT[28]_i_11_n_0 ;
  wire \CRC_OUT[28]_i_3_n_0 ;
  wire \CRC_OUT[28]_i_4_n_0 ;
  wire \CRC_OUT[28]_i_6_n_0 ;
  wire \CRC_OUT[28]_i_7_n_0 ;
  wire \CRC_OUT[2]_i_2_n_0 ;
  wire \CRC_OUT[2]_i_3_n_0 ;
  wire \CRC_OUT[2]_i_4_n_0 ;
  wire \CRC_OUT[2]_i_5_n_0 ;
  wire \CRC_OUT[30]_i_2_n_0 ;
  wire \CRC_OUT[30]_i_3_n_0 ;
  wire \CRC_OUT[30]_i_4_n_0 ;
  wire \CRC_OUT[30]_i_5_n_0 ;
  wire \CRC_OUT[30]_i_6_n_0 ;
  wire \CRC_OUT[30]_i_8_n_0 ;
  wire \CRC_OUT[31]_i_11_n_0 ;
  wire \CRC_OUT[31]_i_3_n_0 ;
  wire \CRC_OUT[31]_i_5_n_0 ;
  wire \CRC_OUT[31]_i_6_n_0 ;
  wire \CRC_OUT[31]_i_7_n_0 ;
  wire \CRC_OUT[31]_i_8_n_0 ;
  wire \CRC_OUT[31]_i_9_n_0 ;
  wire \CRC_OUT[3]_i_2_n_0 ;
  wire \CRC_OUT[3]_i_3_n_0 ;
  wire \CRC_OUT[4]_i_2_n_0 ;
  wire \CRC_OUT[4]_i_3_n_0 ;
  wire \CRC_OUT[4]_i_4_n_0 ;
  wire \CRC_OUT[5]_i_2_n_0 ;
  wire \CRC_OUT[5]_i_4_n_0 ;
  wire \CRC_OUT[5]_i_6_n_0 ;
  wire \CRC_OUT[6]_i_3_n_0 ;
  wire \CRC_OUT[7]_i_2_n_0 ;
  wire \CRC_OUT[7]_i_3_n_0 ;
  wire \CRC_OUT[7]_i_4_n_0 ;
  wire \CRC_OUT[8]_i_2_n_0 ;
  wire \CRC_OUT[8]_i_3_n_0 ;
  wire \CRC_OUT[8]_i_4_n_0 ;
  wire \CRC_OUT[8]_i_5_n_0 ;
  wire \CRC_OUT[9]_i_2_n_0 ;
  wire \CRC_OUT[9]_i_3_n_0 ;
  wire \CRC_OUT[9]_i_4_n_0 ;
  wire \CRC_OUT[9]_i_5_n_0 ;
  wire \CRC_OUT[9]_i_6_n_0 ;
  wire \CRC_OUT_reg[10] ;
  wire \CRC_OUT_reg[11] ;
  wire \CRC_OUT_reg[11]_0 ;
  wire \CRC_OUT_reg[12] ;
  wire \CRC_OUT_reg[13] ;
  wire \CRC_OUT_reg[13]_0 ;
  wire \CRC_OUT_reg[14] ;
  wire \CRC_OUT_reg[14]_0 ;
  wire \CRC_OUT_reg[15] ;
  wire \CRC_OUT_reg[15]_0 ;
  wire \CRC_OUT_reg[16] ;
  wire \CRC_OUT_reg[17] ;
  wire \CRC_OUT_reg[18] ;
  wire \CRC_OUT_reg[18]_0 ;
  wire \CRC_OUT_reg[18]_1 ;
  wire \CRC_OUT_reg[18]_2 ;
  wire [29:0]\CRC_OUT_reg[1] ;
  wire \CRC_OUT_reg[1]_0 ;
  wire \CRC_OUT_reg[20] ;
  wire \CRC_OUT_reg[22] ;
  wire \CRC_OUT_reg[22]_0 ;
  wire \CRC_OUT_reg[23] ;
  wire \CRC_OUT_reg[24] ;
  wire \CRC_OUT_reg[24]_0 ;
  wire \CRC_OUT_reg[25] ;
  wire \CRC_OUT_reg[26] ;
  wire [30:0]\CRC_OUT_reg[27] ;
  wire \CRC_OUT_reg[28] ;
  wire \CRC_OUT_reg[28]_0 ;
  wire \CRC_OUT_reg[30] ;
  wire \CRC_OUT_reg[31] ;
  wire \CRC_OUT_reg[4] ;
  wire \CRC_OUT_reg[5] ;
  wire \CRC_OUT_reg[5]_0 ;
  wire \CRC_OUT_reg[5]_1 ;
  wire \CRC_OUT_reg[6] ;
  wire \CRC_OUT_reg[6]_0 ;
  wire \CRC_OUT_reg[6]_1 ;
  wire \CRC_OUT_reg[8] ;
  wire \CRC_OUT_reg[8]_0 ;
  wire \CRC_OUT_reg[8]_1 ;
  wire \CRC_OUT_reg[8]_2 ;
  wire \CRC_OUT_reg[9] ;
  wire \CRC_OUT_reg[9]_0 ;
  wire \CRC_OUT_reg[9]_1 ;
  wire [5:0]D;
  wire [0:0]E;
  wire [0:0]\FSM_sequential_fifo_state_reg[0]_0 ;
  wire [1:0]Q;
  wire [0:0]SS;
  wire bad_frame_get;
  wire bad_frame_get_reg;
  wire broad_valid_i_10_n_0;
  wire broad_valid_i_2_n_0;
  wire broad_valid_i_3_n_0;
  wire broad_valid_i_4_n_0;
  wire broad_valid_i_5_n_0;
  wire broad_valid_i_6_n_0;
  wire broad_valid_i_7_n_0;
  wire broad_valid_i_8_n_0;
  wire broad_valid_i_9_n_0;
  wire [1:0]\bytes_cnt_reg[1] ;
  wire \bytes_cnt_reg[2] ;
  wire check_reset;
  wire check_reset_i_1_n_0;
  wire check_reset_reg_0;
  wire clk_i;
  wire [47:0]da_addr;
  wire \da_addr_reg[40]_0 ;
  wire \da_addr_reg[6]_0 ;
  wire do_crc_check_reg;
  wire fifo_rd_en;
  wire fifo_rd_en_reg_n_0;
  wire [1:1]fifo_state;
  wire [7:0]get_e_chk;
  wire [7:0]\get_e_chk_reg[7]_0 ;
  wire get_error_code;
  wire get_error_code_i_1_n_0;
  wire get_error_code_i_3_n_0;
  wire get_error_code_reg_0;
  wire get_sfd;
  wire get_sfd0;
  wire get_terminator;
  wire get_terminator_d1;
  wire get_terminator_d2;
  wire get_terminator_d2_reg;
  wire get_terminator_d3;
  wire [0:0]get_terminator_reg_0;
  wire good_frame_get;
  wire good_frame_get_reg;
  wire [0:0]in0;
  wire inband_fcs;
  wire \lt_data_reg_n_0_[10] ;
  wire \lt_data_reg_n_0_[11] ;
  wire \lt_data_reg_n_0_[12] ;
  wire \lt_data_reg_n_0_[13] ;
  wire \lt_data_reg_n_0_[14] ;
  wire \lt_data_reg_n_0_[15] ;
  wire \lt_data_reg_n_0_[1] ;
  wire \lt_data_reg_n_0_[2] ;
  wire \lt_data_reg_n_0_[3] ;
  wire \lt_data_reg_n_0_[4] ;
  wire \lt_data_reg_n_0_[5] ;
  wire \lt_data_reg_n_0_[6] ;
  wire \lt_data_reg_n_0_[7] ;
  wire \lt_data_reg_n_0_[8] ;
  wire \lt_data_reg_n_0_[9] ;
  wire multi_valid_i_10_n_0;
  wire multi_valid_i_2_n_0;
  wire multi_valid_i_3_n_0;
  wire multi_valid_i_4_n_0;
  wire multi_valid_i_5_n_0;
  wire multi_valid_i_6_n_0;
  wire multi_valid_i_7_n_0;
  wire multi_valid_i_8_n_0;
  wire multi_valid_i_9_n_0;
  wire [2:0]pad_cnt;
  wire \pad_cnt[2]_i_2_n_0 ;
  wire [2:0]pad_cnt_reg;
  wire pad_cnt_reg1;
  wire \pad_cnt_reg_n_0_[0] ;
  wire \pad_cnt_reg_n_0_[1] ;
  wire \pad_cnt_reg_n_0_[2] ;
  wire pad_frame;
  wire pad_frame_d1_reg_n_0;
  wire pad_frame_i_2_n_0;
  wire pad_frame_i_3_n_0;
  wire pad_frame_reg_n_0;
  wire [5:3]pad_integer1;
  wire \pad_integer_reg_n_0_[0] ;
  wire \pad_integer_reg_n_0_[1] ;
  wire \pad_integer_reg_n_0_[2] ;
  wire [6:0]pad_last_rxc;
  wire \pad_last_rxc_reg_n_0_[0] ;
  wire \pad_last_rxc_reg_n_0_[1] ;
  wire \pad_last_rxc_reg_n_0_[2] ;
  wire \pad_last_rxc_reg_n_0_[3] ;
  wire \pad_last_rxc_reg_n_0_[4] ;
  wire \pad_last_rxc_reg_n_0_[5] ;
  wire \pad_last_rxc_reg_n_0_[6] ;
  wire [2:0]pad_remain;
  wire [2:0]pad_remain0;
  wire [6:0]pad_rxc_reg;
  wire [71:0]qvDataOut;
  wire receiving;
  wire receiving_d2;
  wire recv_rst;
  wire reset_dcm;
  wire rst_i;
  wire [63:0]\rx_data_reg[63]_0 ;
  wire \rx_data_valid[0]_i_2_n_0 ;
  wire \rx_data_valid[6]_i_2_n_0 ;
  wire \rx_data_valid[6]_i_3_n_0 ;
  wire [7:0]\rx_data_valid_reg[7]_0 ;
  wire [7:0]rxc8_d1;
  wire [7:0]rxc8_d2;
  wire [7:0]rxc8_d3;
  wire [7:0]rxc_end_data;
  wire [7:0]rxc_final;
  wire \rxc_final[0]_i_1_n_0 ;
  wire \rxc_final[1]_i_1_n_0 ;
  wire \rxc_final[2]_i_1_n_0 ;
  wire \rxc_final[3]_i_1_n_0 ;
  wire \rxc_final[4]_i_1_n_0 ;
  wire \rxc_final[5]_i_1_n_0 ;
  wire \rxc_final[6]_i_1_n_0 ;
  wire \rxc_final[7]_i_1_n_0 ;
  wire rxcntrlin_n_0;
  wire rxcntrlin_n_1;
  wire rxcntrlin_n_10;
  wire rxcntrlin_n_2;
  wire rxcntrlin_n_3;
  wire rxcntrlin_n_4;
  wire rxcntrlin_n_5;
  wire rxcntrlin_n_6;
  wire rxcntrlin_n_7;
  wire rxcntrlin_n_8;
  wire rxcntrlin_n_9;
  wire [63:0]rxd64_d1;
  wire [63:0]rxd64_d2;
  wire [63:0]rxd64_d3;
  wire \rxd64_d3_reg[20]_0 ;
  wire \rxd64_d3_reg[29]_0 ;
  wire \rxd64_d3_reg[30]_0 ;
  wire \rxd64_d3_reg[34]_0 ;
  wire \rxd64_d3_reg[40]_0 ;
  wire \rxd64_d3_reg[8]_0 ;
  wire \rxd64_d3_reg[9]_0 ;
  wire rxdatain_n_1;
  wire rxdatain_n_10;
  wire rxdatain_n_11;
  wire rxdatain_n_12;
  wire rxdatain_n_13;
  wire rxdatain_n_14;
  wire rxdatain_n_15;
  wire rxdatain_n_16;
  wire rxdatain_n_17;
  wire rxdatain_n_18;
  wire rxdatain_n_19;
  wire rxdatain_n_2;
  wire rxdatain_n_20;
  wire rxdatain_n_21;
  wire rxdatain_n_22;
  wire rxdatain_n_23;
  wire rxdatain_n_24;
  wire rxdatain_n_25;
  wire rxdatain_n_26;
  wire rxdatain_n_27;
  wire rxdatain_n_28;
  wire rxdatain_n_29;
  wire rxdatain_n_3;
  wire rxdatain_n_30;
  wire rxdatain_n_31;
  wire rxdatain_n_32;
  wire rxdatain_n_33;
  wire rxdatain_n_34;
  wire rxdatain_n_35;
  wire rxdatain_n_36;
  wire rxdatain_n_37;
  wire rxdatain_n_38;
  wire rxdatain_n_39;
  wire rxdatain_n_40;
  wire rxdatain_n_41;
  wire rxdatain_n_42;
  wire rxdatain_n_43;
  wire rxdatain_n_44;
  wire rxdatain_n_45;
  wire rxdatain_n_46;
  wire rxdatain_n_47;
  wire rxdatain_n_48;
  wire rxdatain_n_49;
  wire rxdatain_n_50;
  wire rxdatain_n_51;
  wire rxdatain_n_52;
  wire rxdatain_n_53;
  wire rxdatain_n_54;
  wire rxdatain_n_55;
  wire rxdatain_n_56;
  wire rxdatain_n_57;
  wire rxdatain_n_58;
  wire rxdatain_n_59;
  wire rxdatain_n_6;
  wire rxdatain_n_60;
  wire rxdatain_n_61;
  wire rxdatain_n_62;
  wire rxdatain_n_63;
  wire rxdatain_n_64;
  wire rxdatain_n_65;
  wire rxdatain_n_66;
  wire rxdatain_n_67;
  wire rxdatain_n_68;
  wire rxdatain_n_69;
  wire rxdatain_n_7;
  wire rxdatain_n_70;
  wire rxdatain_n_8;
  wire rxdatain_n_9;
  wire rxfifo_empty;
  wire tagged_frame;
  wire tagged_frame_reg_0;
  wire [1:0]\terminator_location_reg[1]_0 ;
  wire [2:0]\terminator_location_reg[2]_0 ;
  wire [2:0]\terminator_location_reg[2]_1 ;
  wire this_cycle;
  wire this_cycle_reg_n_0;
  wire [7:0]vDataIn;
  wire wait_crc_check;

  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[0]_i_1 
       (.I0(\CRC_OUT[0]_i_2_n_0 ),
        .I1(\CRC_OUT[20]_i_2_n_0 ),
        .I2(\CRC_OUT[12]_i_2_n_0 ),
        .I3(\CRC_OUT[0]_i_3_n_0 ),
        .I4(\CRC_OUT_reg[14] ),
        .I5(\CRC_OUT[0]_i_4_n_0 ),
        .O(\CRC_OUT_reg[27] [0]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[0]_i_2 
       (.I0(\CRC_OUT[10]_i_3_n_0 ),
        .I1(\CRC_OUT[22]_i_6_n_0 ),
        .I2(rxd64_d3[57]),
        .I3(rxd64_d3[63]),
        .I4(\CRC_OUT[31]_i_11_n_0 ),
        .I5(\CRC_OUT_reg[13] ),
        .O(\CRC_OUT[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[0]_i_3 
       (.I0(rxd64_d3[33]),
        .I1(rxd64_d3[35]),
        .O(\CRC_OUT[0]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[0]_i_4 
       (.I0(\CRC_OUT[7]_i_4_n_0 ),
        .I1(rxd64_d3[34]),
        .I2(\CRC_OUT_reg[1] [14]),
        .I3(rxd64_d3[16]),
        .O(\CRC_OUT[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[10]_i_1 
       (.I0(\CRC_OUT[10]_i_2_n_0 ),
        .I1(\CRC_OUT[10]_i_3_n_0 ),
        .I2(\CRC_OUT_reg[10] ),
        .I3(\CRC_OUT[10]_i_5_n_0 ),
        .I4(\CRC_OUT[11]_i_6_n_0 ),
        .I5(\CRC_OUT[27]_i_5_n_0 ),
        .O(\CRC_OUT_reg[27] [10]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[10]_i_2 
       (.I0(\CRC_OUT_reg[1] [23]),
        .I1(rxd64_d3[7]),
        .I2(\rxd64_d3_reg[30]_0 ),
        .I3(rxd64_d3[61]),
        .I4(\CRC_OUT_reg[1] [19]),
        .I5(rxd64_d3[11]),
        .O(\CRC_OUT[10]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[10]_i_3 
       (.I0(rxd64_d3[31]),
        .I1(\CRC_OUT_reg[1] [0]),
        .I2(rxd64_d3[5]),
        .I3(\CRC_OUT_reg[1] [25]),
        .O(\CRC_OUT[10]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[10]_i_5 
       (.I0(rxd64_d3[50]),
        .I1(rxd64_d3[58]),
        .I2(\CRC_OUT_reg[30] ),
        .I3(\CRC_OUT_reg[18] ),
        .I4(\CRC_OUT[26]_i_2_n_0 ),
        .O(\CRC_OUT[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_1 
       (.I0(\CRC_OUT[11]_i_2_n_0 ),
        .I1(\CRC_OUT[11]_i_3_n_0 ),
        .I2(\CRC_OUT[11]_i_4_n_0 ),
        .I3(\CRC_OUT[11]_i_5_n_0 ),
        .I4(\CRC_OUT[11]_i_6_n_0 ),
        .I5(\CRC_OUT_reg[11] ),
        .O(\CRC_OUT_reg[27] [11]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_2 
       (.I0(\CRC_OUT_reg[1] [8]),
        .I1(rxd64_d3[23]),
        .I2(rxd64_d3[20]),
        .I3(\CRC_OUT_reg[1] [10]),
        .I4(rxd64_d3[47]),
        .I5(\rxd64_d3_reg[30]_0 ),
        .O(\CRC_OUT[11]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[11]_i_3 
       (.I0(rxd64_d3[43]),
        .I1(rxd64_d3[59]),
        .O(\CRC_OUT[11]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[11]_i_4 
       (.I0(rxd64_d3[60]),
        .I1(rxd64_d3[35]),
        .O(\CRC_OUT[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[11]_i_5 
       (.I0(\CRC_OUT[28]_i_4_n_0 ),
        .I1(\CRC_OUT_reg[1] [15]),
        .I2(rxd64_d3[15]),
        .I3(\CRC_OUT_reg[11]_0 ),
        .I4(\CRC_OUT[31]_i_3_n_0 ),
        .I5(\CRC_OUT[24]_i_2_n_0 ),
        .O(\CRC_OUT[11]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[11]_i_6 
       (.I0(rxd64_d3[63]),
        .I1(\CRC_OUT[22]_i_5_n_0 ),
        .I2(rxd64_d3[37]),
        .I3(\CRC_OUT_reg[1] [22]),
        .I4(rxd64_d3[8]),
        .O(\CRC_OUT[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[12]_i_1 
       (.I0(\CRC_OUT[20]_i_4_n_0 ),
        .I1(\CRC_OUT[12]_i_2_n_0 ),
        .I2(\CRC_OUT[12]_i_3_n_0 ),
        .I3(\CRC_OUT_reg[12] ),
        .I4(\CRC_OUT[23]_i_5_n_0 ),
        .I5(\CRC_OUT_reg[9] ),
        .O(\CRC_OUT_reg[27] [12]));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[12]_i_2 
       (.I0(rxd64_d3[32]),
        .I1(rxd64_d3[54]),
        .I2(rxd64_d3[0]),
        .I3(\CRC_OUT_reg[1] [29]),
        .O(\CRC_OUT[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[12]_i_3 
       (.I0(\CRC_OUT[31]_i_3_n_0 ),
        .I1(\CRC_OUT_reg[26] ),
        .I2(rxd64_d3[45]),
        .I3(rxd64_d3[61]),
        .I4(rxd64_d3[58]),
        .I5(rxd64_d3[42]),
        .O(\CRC_OUT[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_1 
       (.I0(\CRC_OUT[13]_i_2_n_0 ),
        .I1(\CRC_OUT[13]_i_3_n_0 ),
        .I2(\CRC_OUT[13]_i_4_n_0 ),
        .I3(\CRC_OUT[13]_i_5_n_0 ),
        .I4(\CRC_OUT[30]_i_5_n_0 ),
        .I5(\CRC_OUT[13]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [13]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_2 
       (.I0(\CRC_OUT_reg[10] ),
        .I1(\rxd64_d3_reg[20]_0 ),
        .I2(rxd64_d3[58]),
        .I3(rxd64_d3[38]),
        .I4(\CRC_OUT_reg[13] ),
        .I5(rxd64_d3[53]),
        .O(\CRC_OUT[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[13]_i_3 
       (.I0(rxd64_d3[57]),
        .I1(rxd64_d3[50]),
        .I2(rxd64_d3[45]),
        .I3(rxd64_d3[61]),
        .I4(\CRC_OUT_reg[18] ),
        .I5(\CRC_OUT[11]_i_4_n_0 ),
        .O(\CRC_OUT[13]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[13]_i_4 
       (.I0(rxd64_d3[8]),
        .I1(\CRC_OUT_reg[1] [22]),
        .I2(rxd64_d3[62]),
        .O(\CRC_OUT[13]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[13]_i_5 
       (.I0(rxd64_d3[41]),
        .I1(\CRC_OUT_reg[1] [9]),
        .I2(rxd64_d3[21]),
        .I3(\CRC_OUT_reg[8]_0 ),
        .O(\CRC_OUT[13]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[13]_i_6 
       (.I0(rxd64_d3[32]),
        .I1(rxd64_d3[44]),
        .I2(rxd64_d3[15]),
        .I3(\CRC_OUT_reg[1] [15]),
        .I4(\CRC_OUT_reg[13]_0 ),
        .O(\CRC_OUT[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[14]_i_1 
       (.I0(\CRC_OUT[14]_i_2_n_0 ),
        .I1(\CRC_OUT[19]_i_5_n_0 ),
        .I2(\CRC_OUT[30]_i_5_n_0 ),
        .I3(\CRC_OUT_reg[14] ),
        .I4(\CRC_OUT[14]_i_3_n_0 ),
        .I5(\CRC_OUT[14]_i_4_n_0 ),
        .O(\CRC_OUT_reg[27] [14]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[14]_i_2 
       (.I0(\CRC_OUT[14]_i_5_n_0 ),
        .I1(\CRC_OUT[11]_i_3_n_0 ),
        .I2(\CRC_OUT_reg[17] ),
        .I3(\CRC_OUT[25]_i_8_n_0 ),
        .I4(\CRC_OUT_reg[8]_0 ),
        .I5(\CRC_OUT_reg[14]_0 ),
        .O(\CRC_OUT[14]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[14]_i_3 
       (.I0(rxd64_d3[57]),
        .I1(rxd64_d3[61]),
        .O(\CRC_OUT[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[14]_i_4 
       (.I0(rxd64_d3[52]),
        .I1(\rxd64_d3_reg[20]_0 ),
        .I2(rxd64_d3[40]),
        .I3(rxd64_d3[46]),
        .I4(\CRC_OUT_reg[1] [23]),
        .I5(rxd64_d3[7]),
        .O(\CRC_OUT[14]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[14]_i_5 
       (.I0(rxd64_d3[44]),
        .I1(rxd64_d3[34]),
        .O(\CRC_OUT[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[15]_i_1 
       (.I0(\CRC_OUT[15]_i_2_n_0 ),
        .I1(\CRC_OUT[20]_i_2_n_0 ),
        .I2(\CRC_OUT[15]_i_3_n_0 ),
        .I3(\CRC_OUT[19]_i_5_n_0 ),
        .I4(\CRC_OUT_reg[28]_0 ),
        .O(\CRC_OUT_reg[27] [15]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[15]_i_2 
       (.I0(\CRC_OUT_reg[15] ),
        .I1(\CRC_OUT[15]_i_4_n_0 ),
        .I2(rxd64_d3[45]),
        .I3(rxd64_d3[54]),
        .I4(\CRC_OUT_reg[15]_0 ),
        .I5(rxd64_d3[33]),
        .O(\CRC_OUT[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[15]_i_3 
       (.I0(\CRC_OUT[22]_i_6_n_0 ),
        .I1(\CRC_OUT[27]_i_2_n_0 ),
        .I2(\CRC_OUT_reg[1] [12]),
        .I3(rxd64_d3[18]),
        .I4(\CRC_OUT[27]_i_7_n_0 ),
        .O(\CRC_OUT[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[15]_i_4 
       (.I0(rxd64_d3[6]),
        .I1(\CRC_OUT_reg[1] [24]),
        .O(\CRC_OUT[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[16]_i_1 
       (.I0(\CRC_OUT[16]_i_2_n_0 ),
        .I1(\CRC_OUT[16]_i_3_n_0 ),
        .I2(\CRC_OUT_reg[16] ),
        .I3(rxd64_d3[46]),
        .I4(\CRC_OUT_reg[1] [23]),
        .I5(rxd64_d3[7]),
        .O(\CRC_OUT_reg[27] [16]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[16]_i_2 
       (.I0(\CRC_OUT[16]_i_4_n_0 ),
        .I1(\CRC_OUT[16]_i_5_n_0 ),
        .I2(rxd64_d3[59]),
        .I3(rxd64_d3[41]),
        .I4(rxd64_d3[50]),
        .I5(rxd64_d3[37]),
        .O(\CRC_OUT[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[16]_i_3 
       (.I0(\CRC_OUT[22]_i_4_n_0 ),
        .I1(\CRC_OUT_reg[24]_0 ),
        .I2(\CRC_OUT[28]_i_4_n_0 ),
        .I3(rxd64_d3[33]),
        .I4(rxd64_d3[55]),
        .O(\CRC_OUT[16]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[16]_i_4 
       (.I0(rxd64_d3[58]),
        .I1(rxd64_d3[42]),
        .O(\CRC_OUT[16]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[16]_i_5 
       (.I0(rxd64_d3[17]),
        .I1(\CRC_OUT_reg[1] [13]),
        .I2(rxd64_d3[63]),
        .O(\CRC_OUT[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_1 
       (.I0(\CRC_OUT[17]_i_2_n_0 ),
        .I1(\CRC_OUT[17]_i_3_n_0 ),
        .I2(\CRC_OUT[17]_i_4_n_0 ),
        .I3(\CRC_OUT_reg[16] ),
        .I4(rxd64_d3[43]),
        .I5(rxd64_d3[41]),
        .O(\CRC_OUT_reg[27] [17]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_2 
       (.I0(rxd64_d3[45]),
        .I1(rxd64_d3[33]),
        .I2(rxd64_d3[40]),
        .I3(rxd64_d3[58]),
        .I4(rxd64_d3[36]),
        .I5(rxd64_d3[62]),
        .O(\CRC_OUT[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[17]_i_3 
       (.I0(\CRC_OUT[17]_i_6_n_0 ),
        .I1(\CRC_OUT[22]_i_5_n_0 ),
        .I2(\CRC_OUT_reg[17] ),
        .I3(\CRC_OUT_reg[15]_0 ),
        .I4(\CRC_OUT[26]_i_7_n_0 ),
        .I5(\rxd64_d3_reg[30]_0 ),
        .O(\CRC_OUT[17]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[17]_i_4 
       (.I0(rxd64_d3[38]),
        .I1(\CRC_OUT_reg[1] [12]),
        .I2(rxd64_d3[18]),
        .I3(rxd64_d3[5]),
        .I4(\CRC_OUT_reg[1] [25]),
        .O(\CRC_OUT[17]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_6 
       (.I0(rxd64_d3[57]),
        .I1(rxd64_d3[50]),
        .O(\CRC_OUT[17]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[17]_i_8 
       (.I0(rxd64_d3[30]),
        .I1(\CRC_OUT_reg[1] [1]),
        .O(\rxd64_d3_reg[30]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[18]_i_1 
       (.I0(\CRC_OUT[26]_i_5_n_0 ),
        .I1(\CRC_OUT[18]_i_2_n_0 ),
        .I2(\CRC_OUT[18]_i_3_n_0 ),
        .I3(\CRC_OUT_reg[18]_0 ),
        .I4(\CRC_OUT_reg[18]_1 ),
        .I5(\CRC_OUT[20]_i_5_n_0 ),
        .O(\CRC_OUT_reg[27] [18]));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[18]_i_2 
       (.I0(rxd64_d3[37]),
        .I1(rxd64_d3[39]),
        .O(\CRC_OUT[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[18]_i_3 
       (.I0(\CRC_OUT[14]_i_3_n_0 ),
        .I1(\CRC_OUT[10]_i_3_n_0 ),
        .I2(\CRC_OUT[27]_i_7_n_0 ),
        .I3(rxd64_d3[49]),
        .I4(\CRC_OUT_reg[18]_2 ),
        .I5(\CRC_OUT_reg[5] ),
        .O(\CRC_OUT[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[19]_i_1 
       (.I0(\CRC_OUT[19]_i_2_n_0 ),
        .I1(\CRC_OUT[19]_i_3_n_0 ),
        .I2(\CRC_OUT_reg[18] ),
        .I3(\CRC_OUT[19]_i_5_n_0 ),
        .I4(\CRC_OUT[25]_i_4_n_0 ),
        .I5(\CRC_OUT[19]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [19]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[19]_i_2 
       (.I0(\CRC_OUT[24]_i_8_n_0 ),
        .I1(\CRC_OUT_reg[17] ),
        .I2(rxd64_d3[56]),
        .I3(rxd64_d3[38]),
        .I4(rxd64_d3[36]),
        .I5(rxd64_d3[39]),
        .O(\CRC_OUT[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[19]_i_3 
       (.I0(\CRC_OUT_reg[1] [0]),
        .I1(rxd64_d3[31]),
        .I2(rxd64_d3[28]),
        .I3(\CRC_OUT_reg[1] [3]),
        .I4(rxd64_d3[41]),
        .I5(rxd64_d3[43]),
        .O(\CRC_OUT[19]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[19]_i_4 
       (.I0(\CRC_OUT_reg[1] [17]),
        .I1(rxd64_d3[13]),
        .I2(rxd64_d3[3]),
        .I3(\CRC_OUT_reg[1] [27]),
        .I4(rxd64_d3[47]),
        .O(\CRC_OUT_reg[18] ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[19]_i_5 
       (.I0(rxd64_d3[60]),
        .I1(\CRC_OUT_reg[1] [1]),
        .I2(rxd64_d3[30]),
        .I3(rxd64_d3[55]),
        .I4(\CRC_OUT[31]_i_3_n_0 ),
        .O(\CRC_OUT[19]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[19]_i_6 
       (.I0(rxd64_d3[16]),
        .I1(\CRC_OUT_reg[1] [14]),
        .I2(rxd64_d3[34]),
        .O(\CRC_OUT[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[1]_i_1 
       (.I0(\CRC_OUT[1]_i_2_n_0 ),
        .I1(\CRC_OUT[8]_i_2_n_0 ),
        .I2(\CRC_OUT[1]_i_3_n_0 ),
        .I3(\CRC_OUT_reg[1]_0 ),
        .I4(\CRC_OUT[23]_i_5_n_0 ),
        .I5(\CRC_OUT[28]_i_4_n_0 ),
        .O(\CRC_OUT_reg[27] [1]));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[1]_i_2 
       (.I0(rxd64_d3[1]),
        .I1(\CRC_OUT_reg[1] [28]),
        .I2(rxd64_d3[14]),
        .I3(\CRC_OUT_reg[1] [16]),
        .O(\CRC_OUT[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[1]_i_3 
       (.I0(\CRC_OUT[27]_i_7_n_0 ),
        .I1(\CRC_OUT_reg[18] ),
        .I2(\CRC_OUT_reg[1] [29]),
        .I3(rxd64_d3[0]),
        .I4(rxd64_d3[26]),
        .I5(\CRC_OUT_reg[1] [5]),
        .O(\CRC_OUT[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[20]_i_1 
       (.I0(\CRC_OUT[20]_i_2_n_0 ),
        .I1(\CRC_OUT_reg[14] ),
        .I2(\CRC_OUT_reg[9]_0 ),
        .I3(\CRC_OUT[20]_i_3_n_0 ),
        .I4(\CRC_OUT[20]_i_4_n_0 ),
        .I5(\CRC_OUT[20]_i_5_n_0 ),
        .O(\CRC_OUT_reg[27] [20]));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[20]_i_2 
       (.I0(\CRC_OUT_reg[18] ),
        .I1(rxd64_d3[29]),
        .I2(\CRC_OUT_reg[1] [2]),
        .O(\CRC_OUT[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[20]_i_3 
       (.I0(\CRC_OUT[4]_i_4_n_0 ),
        .I1(\CRC_OUT[0]_i_3_n_0 ),
        .I2(rxd64_d3[46]),
        .I3(rxd64_d3[38]),
        .I4(\CRC_OUT_reg[20] ),
        .I5(rxd64_d3[54]),
        .O(\CRC_OUT[20]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[20]_i_4 
       (.I0(rxd64_d3[59]),
        .I1(rxd64_d3[51]),
        .O(\CRC_OUT[20]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[20]_i_5 
       (.I0(rxd64_d3[40]),
        .I1(rxd64_d3[42]),
        .O(\CRC_OUT[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[21]_i_1 
       (.I0(\CRC_OUT_reg[28]_0 ),
        .I1(\CRC_OUT[30]_i_4_n_0 ),
        .I2(\CRC_OUT[21]_i_2_n_0 ),
        .I3(rxd64_d3[39]),
        .I4(rxd64_d3[37]),
        .I5(\CRC_OUT[21]_i_3_n_0 ),
        .O(\CRC_OUT_reg[27] [21]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[21]_i_2 
       (.I0(\CRC_OUT_reg[9] ),
        .I1(\CRC_OUT[21]_i_4_n_0 ),
        .I2(\rxd64_d3_reg[29]_0 ),
        .I3(rxd64_d3[53]),
        .I4(rxd64_d3[26]),
        .I5(\CRC_OUT_reg[1] [5]),
        .O(\CRC_OUT[21]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[21]_i_3 
       (.I0(rxd64_d3[50]),
        .I1(rxd64_d3[58]),
        .O(\CRC_OUT[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[21]_i_4 
       (.I0(\CRC_OUT_reg[1] [8]),
        .I1(rxd64_d3[23]),
        .I2(rxd64_d3[54]),
        .I3(rxd64_d3[32]),
        .I4(rxd64_d3[46]),
        .I5(rxd64_d3[45]),
        .O(\CRC_OUT[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[22]_i_1 
       (.I0(\CRC_OUT[22]_i_2_n_0 ),
        .I1(\CRC_OUT[30]_i_6_n_0 ),
        .I2(\CRC_OUT_reg[22] ),
        .I3(\CRC_OUT[22]_i_4_n_0 ),
        .I4(rxd64_d3[63]),
        .I5(\CRC_OUT[22]_i_5_n_0 ),
        .O(\CRC_OUT_reg[27] [22]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[22]_i_2 
       (.I0(\CRC_OUT_reg[10] ),
        .I1(\CRC_OUT[22]_i_6_n_0 ),
        .I2(rxd64_d3[36]),
        .I3(rxd64_d3[47]),
        .I4(\CRC_OUT_reg[22]_0 ),
        .I5(rxd64_d3[45]),
        .O(\CRC_OUT[22]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[22]_i_4 
       (.I0(rxd64_d3[34]),
        .I1(rxd64_d3[44]),
        .I2(\CRC_OUT_reg[1] [5]),
        .I3(rxd64_d3[26]),
        .O(\CRC_OUT[22]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[22]_i_5 
       (.I0(\CRC_OUT_reg[1] [4]),
        .I1(rxd64_d3[27]),
        .I2(rxd64_d3[54]),
        .I3(rxd64_d3[32]),
        .I4(rxd64_d3[49]),
        .O(\CRC_OUT[22]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[22]_i_6 
       (.I0(rxd64_d3[39]),
        .I1(rxd64_d3[19]),
        .I2(\CRC_OUT_reg[1] [11]),
        .I3(rxd64_d3[51]),
        .O(\CRC_OUT[22]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[22]_i_7 
       (.I0(\CRC_OUT_reg[1] [6]),
        .I1(rxd64_d3[25]),
        .I2(rxd64_d3[52]),
        .O(\CRC_OUT_reg[6] ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[23]_i_1 
       (.I0(\CRC_OUT[23]_i_2_n_0 ),
        .I1(\CRC_OUT[31]_i_3_n_0 ),
        .I2(\rxd64_d3_reg[29]_0 ),
        .I3(\CRC_OUT[23]_i_4_n_0 ),
        .I4(\CRC_OUT[23]_i_5_n_0 ),
        .I5(\CRC_OUT[23]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [23]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[23]_i_2 
       (.I0(\rxd64_d3_reg[8]_0 ),
        .I1(\CRC_OUT_reg[18] ),
        .I2(\CRC_OUT_reg[23] ),
        .I3(rxd64_d3[43]),
        .I4(\CRC_OUT_reg[20] ),
        .I5(\CRC_OUT[26]_i_7_n_0 ),
        .O(\CRC_OUT[23]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[23]_i_3 
       (.I0(rxd64_d3[29]),
        .I1(\CRC_OUT_reg[1] [2]),
        .I2(\CRC_OUT_reg[1] [3]),
        .I3(rxd64_d3[28]),
        .O(\rxd64_d3_reg[29]_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[23]_i_4 
       (.I0(\CRC_OUT_reg[1] [4]),
        .I1(rxd64_d3[27]),
        .I2(rxd64_d3[54]),
        .I3(rxd64_d3[32]),
        .I4(\CRC_OUT[1]_i_2_n_0 ),
        .O(\CRC_OUT[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[23]_i_5 
       (.I0(rxd64_d3[57]),
        .I1(rxd64_d3[50]),
        .I2(rxd64_d3[17]),
        .I3(\CRC_OUT_reg[1] [13]),
        .I4(rxd64_d3[63]),
        .I5(\CRC_OUT[24]_i_2_n_0 ),
        .O(\CRC_OUT[23]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[23]_i_6 
       (.I0(rxd64_d3[34]),
        .I1(rxd64_d3[44]),
        .I2(rxd64_d3[21]),
        .I3(\CRC_OUT_reg[1] [9]),
        .O(\CRC_OUT[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_1 
       (.I0(\CRC_OUT[24]_i_2_n_0 ),
        .I1(\CRC_OUT[24]_i_3_n_0 ),
        .I2(\CRC_OUT[24]_i_4_n_0 ),
        .I3(\CRC_OUT_reg[24] ),
        .I4(\CRC_OUT[24]_i_6_n_0 ),
        .I5(\CRC_OUT_reg[24]_0 ),
        .O(\CRC_OUT_reg[27] [24]));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[24]_i_10 
       (.I0(\CRC_OUT_reg[1] [5]),
        .I1(rxd64_d3[26]),
        .I2(rxd64_d3[53]),
        .O(\CRC_OUT_reg[5] ));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_12 
       (.I0(rxd64_d3[20]),
        .I1(\CRC_OUT_reg[1] [10]),
        .O(\rxd64_d3_reg[20]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[24]_i_2 
       (.I0(rxd64_d3[62]),
        .I1(rxd64_d3[46]),
        .I2(rxd64_d3[36]),
        .I3(\CRC_OUT_reg[1] [23]),
        .I4(rxd64_d3[7]),
        .O(\CRC_OUT[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_3 
       (.I0(\CRC_OUT_reg[1] [8]),
        .I1(rxd64_d3[23]),
        .I2(\CRC_OUT_reg[1] [29]),
        .I3(rxd64_d3[0]),
        .I4(rxd64_d3[35]),
        .I5(rxd64_d3[33]),
        .O(\CRC_OUT[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[24]_i_4 
       (.I0(\CRC_OUT[24]_i_8_n_0 ),
        .I1(\CRC_OUT_reg[15] ),
        .I2(rxd64_d3[56]),
        .I3(rxd64_d3[42]),
        .I4(rxd64_d3[43]),
        .I5(rxd64_d3[49]),
        .O(\CRC_OUT[24]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[24]_i_6 
       (.I0(rxd64_d3[61]),
        .I1(rxd64_d3[45]),
        .I2(rxd64_d3[24]),
        .I3(\CRC_OUT_reg[1] [7]),
        .O(\CRC_OUT[24]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[24]_i_8 
       (.I0(rxd64_d3[12]),
        .I1(\CRC_OUT_reg[1] [18]),
        .O(\CRC_OUT[24]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_1 
       (.I0(\CRC_OUT[25]_i_2_n_0 ),
        .I1(\CRC_OUT[25]_i_3_n_0 ),
        .I2(\CRC_OUT[25]_i_4_n_0 ),
        .I3(\CRC_OUT_reg[9]_0 ),
        .I4(\CRC_OUT[25]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [25]));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_10 
       (.I0(rxd64_d3[45]),
        .I1(rxd64_d3[61]),
        .O(\CRC_OUT[25]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[25]_i_2 
       (.I0(\CRC_OUT_reg[22]_0 ),
        .I1(\CRC_OUT[25]_i_8_n_0 ),
        .I2(rxd64_d3[42]),
        .I3(rxd64_d3[41]),
        .I4(rxd64_d3[32]),
        .I5(rxd64_d3[48]),
        .O(\CRC_OUT[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[25]_i_3 
       (.I0(\CRC_OUT[22]_i_4_n_0 ),
        .I1(\CRC_OUT[25]_i_9_n_0 ),
        .I2(\CRC_OUT_reg[25] ),
        .I3(\CRC_OUT[11]_i_4_n_0 ),
        .I4(\CRC_OUT[25]_i_10_n_0 ),
        .I5(\CRC_OUT[1]_i_2_n_0 ),
        .O(\CRC_OUT[25]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_4 
       (.I0(rxd64_d3[52]),
        .I1(rxd64_d3[25]),
        .I2(\CRC_OUT_reg[1] [6]),
        .I3(rxd64_d3[23]),
        .I4(\CRC_OUT_reg[1] [8]),
        .O(\CRC_OUT[25]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[25]_i_6 
       (.I0(rxd64_d3[55]),
        .I1(rxd64_d3[30]),
        .I2(\CRC_OUT_reg[1] [1]),
        .I3(\CRC_OUT_reg[1] [24]),
        .I4(rxd64_d3[6]),
        .O(\CRC_OUT[25]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[25]_i_8 
       (.I0(rxd64_d3[19]),
        .I1(\CRC_OUT_reg[1] [11]),
        .O(\CRC_OUT[25]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[25]_i_9 
       (.I0(rxd64_d3[7]),
        .I1(\CRC_OUT_reg[1] [23]),
        .I2(rxd64_d3[46]),
        .O(\CRC_OUT[25]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_1 
       (.I0(\CRC_OUT[26]_i_2_n_0 ),
        .I1(\CRC_OUT_reg[26] ),
        .I2(\CRC_OUT_reg[14] ),
        .I3(\CRC_OUT[26]_i_4_n_0 ),
        .I4(\CRC_OUT_reg[31] ),
        .I5(\CRC_OUT[26]_i_5_n_0 ),
        .O(\CRC_OUT_reg[27] [26]));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[26]_i_2 
       (.I0(rxd64_d3[35]),
        .I1(rxd64_d3[60]),
        .I2(rxd64_d3[24]),
        .I3(\CRC_OUT_reg[1] [7]),
        .O(\CRC_OUT[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_4 
       (.I0(\CRC_OUT[26]_i_6_n_0 ),
        .I1(\CRC_OUT[28]_i_11_n_0 ),
        .I2(\CRC_OUT[1]_i_2_n_0 ),
        .I3(\CRC_OUT[26]_i_7_n_0 ),
        .I4(\CRC_OUT[5]_i_4_n_0 ),
        .I5(\CRC_OUT[26]_i_8_n_0 ),
        .O(\CRC_OUT[26]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[26]_i_5 
       (.I0(rxd64_d3[44]),
        .I1(rxd64_d3[32]),
        .O(\CRC_OUT[26]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[26]_i_6 
       (.I0(rxd64_d3[45]),
        .I1(rxd64_d3[57]),
        .I2(rxd64_d3[63]),
        .I3(rxd64_d3[38]),
        .I4(rxd64_d3[53]),
        .I5(rxd64_d3[40]),
        .O(\CRC_OUT[26]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[26]_i_7 
       (.I0(rxd64_d3[25]),
        .I1(\CRC_OUT_reg[1] [6]),
        .O(\CRC_OUT[26]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[26]_i_8 
       (.I0(rxd64_d3[41]),
        .I1(\CRC_OUT_reg[1] [9]),
        .I2(rxd64_d3[21]),
        .I3(rxd64_d3[59]),
        .I4(rxd64_d3[43]),
        .O(\CRC_OUT[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_1 
       (.I0(\CRC_OUT[27]_i_2_n_0 ),
        .I1(\CRC_OUT_reg[14] ),
        .I2(\CRC_OUT[31]_i_7_n_0 ),
        .I3(\CRC_OUT[27]_i_4_n_0 ),
        .I4(\CRC_OUT_reg[28]_0 ),
        .I5(\CRC_OUT[27]_i_5_n_0 ),
        .O(\CRC_OUT_reg[27] [27]));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[27]_i_2 
       (.I0(rxd64_d3[42]),
        .I1(rxd64_d3[58]),
        .I2(rxd64_d3[59]),
        .I3(rxd64_d3[43]),
        .O(\CRC_OUT[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_4 
       (.I0(\CRC_OUT[27]_i_6_n_0 ),
        .I1(\CRC_OUT[27]_i_7_n_0 ),
        .I2(\CRC_OUT[10]_i_3_n_0 ),
        .I3(rxd64_d3[62]),
        .I4(rxd64_d3[39]),
        .I5(\CRC_OUT[27]_i_8_n_0 ),
        .O(\CRC_OUT[27]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[27]_i_5 
       (.I0(\CRC_OUT_reg[1] [9]),
        .I1(rxd64_d3[21]),
        .I2(rxd64_d3[44]),
        .I3(rxd64_d3[34]),
        .I4(\CRC_OUT[28]_i_10_n_0 ),
        .O(\CRC_OUT[27]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[27]_i_6 
       (.I0(rxd64_d3[18]),
        .I1(\CRC_OUT_reg[1] [12]),
        .I2(rxd64_d3[38]),
        .O(\CRC_OUT[27]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[27]_i_7 
       (.I0(\CRC_OUT_reg[1] [20]),
        .I1(rxd64_d3[10]),
        .I2(rxd64_d3[56]),
        .O(\CRC_OUT[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[27]_i_8 
       (.I0(rxd64_d3[24]),
        .I1(\CRC_OUT_reg[1] [7]),
        .I2(\CRC_OUT_reg[1] [17]),
        .I3(rxd64_d3[13]),
        .I4(rxd64_d3[3]),
        .I5(\CRC_OUT_reg[1] [27]),
        .O(\CRC_OUT[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_1 
       (.I0(\CRC_OUT_reg[28] ),
        .I1(\CRC_OUT[28]_i_3_n_0 ),
        .I2(\CRC_OUT[28]_i_4_n_0 ),
        .I3(\CRC_OUT_reg[28]_0 ),
        .I4(\CRC_OUT[28]_i_6_n_0 ),
        .I5(\CRC_OUT[28]_i_7_n_0 ),
        .O(\CRC_OUT_reg[27] [28]));
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_10 
       (.I0(rxd64_d3[0]),
        .I1(\CRC_OUT_reg[1] [29]),
        .I2(rxd64_d3[23]),
        .I3(\CRC_OUT_reg[1] [8]),
        .O(\CRC_OUT[28]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[28]_i_11 
       (.I0(rxd64_d3[9]),
        .I1(\CRC_OUT_reg[1] [21]),
        .I2(rxd64_d3[4]),
        .I3(\CRC_OUT_reg[1] [26]),
        .O(\CRC_OUT[28]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_3 
       (.I0(\CRC_OUT[28]_i_10_n_0 ),
        .I1(rxd64_d3[57]),
        .I2(rxd64_d3[61]),
        .I3(\CRC_OUT[28]_i_11_n_0 ),
        .I4(rxd64_d3[58]),
        .I5(rxd64_d3[42]),
        .O(\CRC_OUT[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[28]_i_4 
       (.I0(rxd64_d3[51]),
        .I1(\CRC_OUT_reg[1] [11]),
        .I2(rxd64_d3[19]),
        .I3(rxd64_d3[39]),
        .I4(\CRC_OUT_reg[1] [18]),
        .I5(rxd64_d3[12]),
        .O(\CRC_OUT[28]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[28]_i_6 
       (.I0(rxd64_d3[43]),
        .I1(rxd64_d3[41]),
        .O(\CRC_OUT[28]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[28]_i_7 
       (.I0(\CRC_OUT_reg[1] [13]),
        .I1(rxd64_d3[17]),
        .I2(rxd64_d3[33]),
        .I3(rxd64_d3[35]),
        .I4(\CRC_OUT[25]_i_6_n_0 ),
        .O(\CRC_OUT[28]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[29]_i_3 
       (.I0(rxd64_d3[8]),
        .I1(\CRC_OUT_reg[1] [22]),
        .I2(rxd64_d3[37]),
        .O(\rxd64_d3_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_5 
       (.I0(rxd64_d3[40]),
        .I1(rxd64_d3[42]),
        .I2(\CRC_OUT[12]_i_2_n_0 ),
        .I3(\CRC_OUT[11]_i_4_n_0 ),
        .I4(rxd64_d3[57]),
        .I5(rxd64_d3[50]),
        .O(\rxd64_d3_reg[40]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[29]_i_6 
       (.I0(rxd64_d3[34]),
        .I1(rxd64_d3[41]),
        .I2(\CRC_OUT_reg[1] [9]),
        .I3(rxd64_d3[21]),
        .I4(\CRC_OUT_reg[8]_0 ),
        .I5(rxd64_d3[56]),
        .O(\rxd64_d3_reg[34]_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[2]_i_1 
       (.I0(\CRC_OUT[2]_i_2_n_0 ),
        .I1(\CRC_OUT[11]_i_6_n_0 ),
        .I2(\CRC_OUT[2]_i_3_n_0 ),
        .O(\CRC_OUT_reg[27] [2]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[2]_i_2 
       (.I0(\CRC_OUT_reg[8]_0 ),
        .I1(\CRC_OUT[5]_i_4_n_0 ),
        .I2(\CRC_OUT[15]_i_4_n_0 ),
        .I3(rxd64_d3[47]),
        .I4(\CRC_OUT[2]_i_4_n_0 ),
        .I5(\CRC_OUT[26]_i_7_n_0 ),
        .O(\CRC_OUT[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[2]_i_3 
       (.I0(\CRC_OUT[2]_i_5_n_0 ),
        .I1(\CRC_OUT[8]_i_5_n_0 ),
        .I2(\CRC_OUT[17]_i_6_n_0 ),
        .I3(\CRC_OUT[24]_i_6_n_0 ),
        .I4(\CRC_OUT[10]_i_3_n_0 ),
        .I5(\CRC_OUT[27]_i_7_n_0 ),
        .O(\CRC_OUT[2]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[2]_i_4 
       (.I0(rxd64_d3[26]),
        .I1(\CRC_OUT_reg[1] [5]),
        .O(\CRC_OUT[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[2]_i_5 
       (.I0(\CRC_OUT_reg[1] [26]),
        .I1(rxd64_d3[4]),
        .I2(rxd64_d3[28]),
        .I3(\CRC_OUT_reg[1] [3]),
        .I4(rxd64_d3[55]),
        .I5(rxd64_d3[33]),
        .O(\CRC_OUT[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[30]_i_1 
       (.I0(\CRC_OUT[30]_i_2_n_0 ),
        .I1(\CRC_OUT[30]_i_3_n_0 ),
        .I2(\CRC_OUT[30]_i_4_n_0 ),
        .I3(\CRC_OUT[30]_i_5_n_0 ),
        .I4(\CRC_OUT[30]_i_6_n_0 ),
        .I5(\CRC_OUT_reg[30] ),
        .O(\CRC_OUT_reg[27] [29]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[30]_i_2 
       (.I0(\CRC_OUT[30]_i_8_n_0 ),
        .I1(\CRC_OUT_reg[25] ),
        .I2(rxd64_d3[53]),
        .I3(rxd64_d3[55]),
        .I4(\CRC_OUT_reg[14]_0 ),
        .I5(rxd64_d3[59]),
        .O(\CRC_OUT[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[30]_i_3 
       (.I0(\CRC_OUT_reg[1] [13]),
        .I1(rxd64_d3[17]),
        .I2(rxd64_d3[33]),
        .I3(rxd64_d3[35]),
        .I4(rxd64_d3[39]),
        .I5(rxd64_d3[37]),
        .O(\CRC_OUT[30]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[30]_i_4 
       (.I0(\CRC_OUT_reg[8]_0 ),
        .I1(rxd64_d3[21]),
        .I2(\CRC_OUT_reg[1] [9]),
        .I3(rxd64_d3[41]),
        .I4(rxd64_d3[34]),
        .O(\CRC_OUT[30]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[30]_i_5 
       (.I0(\CRC_OUT[10]_i_3_n_0 ),
        .I1(\CRC_OUT_reg[1] [20]),
        .I2(rxd64_d3[10]),
        .I3(rxd64_d3[56]),
        .I4(rxd64_d3[49]),
        .O(\CRC_OUT[30]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[30]_i_6 
       (.I0(rxd64_d3[40]),
        .I1(rxd64_d3[20]),
        .I2(\CRC_OUT_reg[1] [10]),
        .I3(rxd64_d3[18]),
        .I4(\CRC_OUT_reg[1] [12]),
        .O(\CRC_OUT[30]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[30]_i_8 
       (.I0(rxd64_d3[7]),
        .I1(\CRC_OUT_reg[1] [23]),
        .I2(rxd64_d3[36]),
        .O(\CRC_OUT[30]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[31]_i_11 
       (.I0(rxd64_d3[10]),
        .I1(\CRC_OUT_reg[1] [20]),
        .O(\CRC_OUT[31]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \CRC_OUT[31]_i_1__2 
       (.I0(get_error_code),
        .I1(get_terminator_d3),
        .I2(rst_i),
        .I3(recv_rst),
        .O(SS));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[31]_i_2 
       (.I0(\CRC_OUT[31]_i_3_n_0 ),
        .I1(\CRC_OUT_reg[31] ),
        .I2(\CRC_OUT[31]_i_5_n_0 ),
        .I3(\CRC_OUT[31]_i_6_n_0 ),
        .I4(\CRC_OUT[31]_i_7_n_0 ),
        .I5(\CRC_OUT[31]_i_8_n_0 ),
        .O(\CRC_OUT_reg[27] [30]));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[31]_i_3 
       (.I0(\CRC_OUT_reg[1] [26]),
        .I1(rxd64_d3[4]),
        .I2(\CRC_OUT_reg[1] [21]),
        .I3(rxd64_d3[9]),
        .I4(rxd64_d3[48]),
        .O(\CRC_OUT[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[31]_i_5 
       (.I0(\CRC_OUT[1]_i_2_n_0 ),
        .I1(\CRC_OUT[31]_i_9_n_0 ),
        .I2(\CRC_OUT_reg[13]_0 ),
        .I3(\CRC_OUT_reg[1] [1]),
        .I4(rxd64_d3[30]),
        .I5(rxd64_d3[55]),
        .O(\CRC_OUT[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[31]_i_6 
       (.I0(\CRC_OUT[31]_i_11_n_0 ),
        .I1(\CRC_OUT[5]_i_4_n_0 ),
        .I2(rxd64_d3[34]),
        .I3(rxd64_d3[38]),
        .I4(rxd64_d3[36]),
        .I5(rxd64_d3[58]),
        .O(\CRC_OUT[31]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_7 
       (.I0(rxd64_d3[40]),
        .I1(rxd64_d3[20]),
        .I2(\CRC_OUT_reg[1] [10]),
        .I3(rxd64_d3[52]),
        .O(\CRC_OUT[31]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_8 
       (.I0(rxd64_d3[35]),
        .I1(rxd64_d3[33]),
        .I2(rxd64_d3[17]),
        .I3(\CRC_OUT_reg[1] [13]),
        .O(\CRC_OUT[31]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[31]_i_9 
       (.I0(rxd64_d3[32]),
        .I1(rxd64_d3[54]),
        .I2(rxd64_d3[27]),
        .I3(\CRC_OUT_reg[1] [4]),
        .O(\CRC_OUT[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[3]_i_1 
       (.I0(\CRC_OUT[7]_i_4_n_0 ),
        .I1(\CRC_OUT[3]_i_2_n_0 ),
        .I2(\CRC_OUT[3]_i_3_n_0 ),
        .I3(\CRC_OUT[24]_i_6_n_0 ),
        .I4(\CRC_OUT[19]_i_5_n_0 ),
        .I5(\CRC_OUT_reg[31] ),
        .O(\CRC_OUT_reg[27] [3]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[3]_i_2 
       (.I0(\CRC_OUT_reg[1] [8]),
        .I1(rxd64_d3[23]),
        .I2(\CRC_OUT[27]_i_7_n_0 ),
        .I3(\CRC_OUT[10]_i_3_n_0 ),
        .I4(rxd64_d3[44]),
        .I5(\CRC_OUT[26]_i_7_n_0 ),
        .O(\CRC_OUT[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[3]_i_3 
       (.I0(rxd64_d3[49]),
        .I1(rxd64_d3[32]),
        .I2(rxd64_d3[54]),
        .I3(rxd64_d3[27]),
        .I4(\CRC_OUT_reg[1] [4]),
        .I5(\CRC_OUT[24]_i_2_n_0 ),
        .O(\CRC_OUT[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_1 
       (.I0(\CRC_OUT[4]_i_2_n_0 ),
        .I1(\CRC_OUT[4]_i_3_n_0 ),
        .I2(\CRC_OUT[4]_i_4_n_0 ),
        .I3(rxd64_d3[60]),
        .I4(\CRC_OUT_reg[11] ),
        .I5(\CRC_OUT_reg[18]_1 ),
        .O(\CRC_OUT_reg[27] [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_2 
       (.I0(\CRC_OUT_reg[4] ),
        .I1(\CRC_OUT[14]_i_5_n_0 ),
        .I2(rxd64_d3[32]),
        .I3(rxd64_d3[48]),
        .I4(rxd64_d3[33]),
        .I5(rxd64_d3[57]),
        .O(\CRC_OUT[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[4]_i_3 
       (.I0(\CRC_OUT[28]_i_10_n_0 ),
        .I1(\CRC_OUT[24]_i_6_n_0 ),
        .I2(\CRC_OUT[11]_i_3_n_0 ),
        .I3(\CRC_OUT[22]_i_6_n_0 ),
        .I4(\CRC_OUT[16]_i_5_n_0 ),
        .I5(\CRC_OUT_reg[6] ),
        .O(\CRC_OUT[4]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[4]_i_4 
       (.I0(\CRC_OUT_reg[1] [1]),
        .I1(rxd64_d3[30]),
        .I2(rxd64_d3[55]),
        .O(\CRC_OUT[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[5]_i_1 
       (.I0(\CRC_OUT[5]_i_2_n_0 ),
        .I1(\CRC_OUT_reg[5]_0 ),
        .I2(\CRC_OUT[5]_i_4_n_0 ),
        .I3(\CRC_OUT_reg[5]_1 ),
        .I4(\CRC_OUT[27]_i_5_n_0 ),
        .I5(\CRC_OUT[5]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[5]_i_2 
       (.I0(\CRC_OUT[26]_i_2_n_0 ),
        .I1(\CRC_OUT[13]_i_4_n_0 ),
        .I2(\CRC_OUT[27]_i_7_n_0 ),
        .I3(\CRC_OUT[28]_i_11_n_0 ),
        .I4(\CRC_OUT[27]_i_2_n_0 ),
        .I5(\CRC_OUT_reg[5] ),
        .O(\CRC_OUT[5]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[5]_i_4 
       (.I0(\CRC_OUT_reg[1] [11]),
        .I1(rxd64_d3[19]),
        .I2(rxd64_d3[39]),
        .O(\CRC_OUT[5]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[5]_i_6 
       (.I0(rxd64_d3[63]),
        .I1(\CRC_OUT_reg[1] [13]),
        .I2(rxd64_d3[17]),
        .I3(rxd64_d3[50]),
        .I4(rxd64_d3[57]),
        .O(\CRC_OUT[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[6]_i_1 
       (.I0(\CRC_OUT_reg[6]_0 ),
        .I1(\CRC_OUT[6]_i_3_n_0 ),
        .I2(rxd64_d3[33]),
        .I3(rxd64_d3[55]),
        .I4(\rxd64_d3_reg[34]_0 ),
        .I5(\CRC_OUT[25]_i_4_n_0 ),
        .O(\CRC_OUT_reg[27] [6]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[6]_i_3 
       (.I0(\CRC_OUT[27]_i_2_n_0 ),
        .I1(\CRC_OUT[13]_i_4_n_0 ),
        .I2(\CRC_OUT_reg[6]_1 ),
        .I3(rxd64_d3[61]),
        .I4(rxd64_d3[57]),
        .I5(\CRC_OUT[27]_i_6_n_0 ),
        .O(\CRC_OUT[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[7]_i_1 
       (.I0(\CRC_OUT[7]_i_2_n_0 ),
        .I1(\CRC_OUT[7]_i_3_n_0 ),
        .I2(\CRC_OUT[20]_i_2_n_0 ),
        .I3(\rxd64_d3_reg[34]_0 ),
        .I4(\CRC_OUT[7]_i_4_n_0 ),
        .O(\CRC_OUT_reg[27] [7]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \CRC_OUT[7]_i_2 
       (.I0(\rxd64_d3_reg[9]_0 ),
        .I1(rxd64_d3[55]),
        .I2(rxd64_d3[61]),
        .I3(rxd64_d3[39]),
        .I4(rxd64_d3[48]),
        .O(\CRC_OUT[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[7]_i_3 
       (.I0(\CRC_OUT_reg[26] ),
        .I1(\CRC_OUT[26]_i_2_n_0 ),
        .I2(\CRC_OUT[16]_i_4_n_0 ),
        .I3(\CRC_OUT[10]_i_3_n_0 ),
        .I4(\CRC_OUT[16]_i_5_n_0 ),
        .I5(\CRC_OUT[9]_i_6_n_0 ),
        .O(\CRC_OUT[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[7]_i_4 
       (.I0(rxd64_d3[53]),
        .I1(rxd64_d3[26]),
        .I2(\CRC_OUT_reg[1] [5]),
        .I3(rxd64_d3[38]),
        .I4(\CRC_OUT_reg[1] [12]),
        .I5(rxd64_d3[18]),
        .O(\CRC_OUT[7]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CRC_OUT[7]_i_5 
       (.I0(rxd64_d3[9]),
        .I1(\CRC_OUT_reg[1] [21]),
        .I2(rxd64_d3[7]),
        .I3(\CRC_OUT_reg[1] [23]),
        .O(\rxd64_d3_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_1 
       (.I0(\CRC_OUT[8]_i_2_n_0 ),
        .I1(\CRC_OUT[20]_i_4_n_0 ),
        .I2(\CRC_OUT[8]_i_3_n_0 ),
        .I3(\CRC_OUT[8]_i_4_n_0 ),
        .I4(\CRC_OUT[25]_i_6_n_0 ),
        .I5(\CRC_OUT[30]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [8]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_2 
       (.I0(rxd64_d3[28]),
        .I1(\CRC_OUT_reg[1] [3]),
        .I2(\CRC_OUT_reg[1] [2]),
        .I3(rxd64_d3[29]),
        .I4(rxd64_d3[52]),
        .I5(\CRC_OUT[26]_i_7_n_0 ),
        .O(\CRC_OUT[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_3 
       (.I0(\CRC_OUT[28]_i_10_n_0 ),
        .I1(rxd64_d3[41]),
        .I2(\CRC_OUT_reg[8] ),
        .I3(\CRC_OUT_reg[8]_0 ),
        .I4(\CRC_OUT_reg[5] ),
        .I5(\CRC_OUT[16]_i_5_n_0 ),
        .O(\CRC_OUT[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[8]_i_4 
       (.I0(\CRC_OUT[11]_i_4_n_0 ),
        .I1(\CRC_OUT[8]_i_5_n_0 ),
        .I2(\CRC_OUT_reg[8]_1 ),
        .I3(rxd64_d3[32]),
        .I4(\CRC_OUT[28]_i_11_n_0 ),
        .I5(\CRC_OUT_reg[8]_2 ),
        .O(\CRC_OUT[8]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[8]_i_5 
       (.I0(rxd64_d3[46]),
        .I1(rxd64_d3[62]),
        .O(\CRC_OUT[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_1 
       (.I0(\CRC_OUT[9]_i_2_n_0 ),
        .I1(\CRC_OUT[9]_i_3_n_0 ),
        .I2(\CRC_OUT[9]_i_4_n_0 ),
        .I3(\CRC_OUT_reg[9] ),
        .I4(\CRC_OUT_reg[9]_0 ),
        .I5(\CRC_OUT[19]_i_6_n_0 ),
        .O(\CRC_OUT_reg[27] [9]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_2 
       (.I0(\CRC_OUT_reg[9]_1 ),
        .I1(\CRC_OUT[10]_i_3_n_0 ),
        .I2(rxd64_d3[54]),
        .I3(rxd64_d3[59]),
        .I4(\rxd64_d3_reg[30]_0 ),
        .I5(\CRC_OUT[9]_i_5_n_0 ),
        .O(\CRC_OUT[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_3 
       (.I0(\CRC_OUT[24]_i_6_n_0 ),
        .I1(rxd64_d3[8]),
        .I2(\CRC_OUT_reg[1] [22]),
        .I3(rxd64_d3[62]),
        .I4(\CRC_OUT[22]_i_6_n_0 ),
        .I5(\CRC_OUT[9]_i_6_n_0 ),
        .O(\CRC_OUT[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CRC_OUT[9]_i_4 
       (.I0(rxd64_d3[58]),
        .I1(rxd64_d3[50]),
        .I2(\CRC_OUT_reg[1] [6]),
        .I3(rxd64_d3[25]),
        .I4(rxd64_d3[52]),
        .I5(\rxd64_d3_reg[29]_0 ),
        .O(\CRC_OUT[9]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CRC_OUT[9]_i_5 
       (.I0(rxd64_d3[3]),
        .I1(\CRC_OUT_reg[1] [27]),
        .O(\CRC_OUT[9]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CRC_OUT[9]_i_6 
       (.I0(\CRC_OUT_reg[1] [10]),
        .I1(rxd64_d3[20]),
        .I2(rxd64_d3[40]),
        .O(\CRC_OUT[9]_i_6_n_0 ));
  (* FSM_ENCODED_STATES = "WAIT_TMP:10,READ:11,IDLE:01,WAIT:00" *) 
  FDPE #(
    .INIT(1'b1)) 
    \FSM_sequential_fifo_state_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(rxcntrlin_n_1),
        .PRE(reset_dcm),
        .Q(\FSM_sequential_fifo_state_reg[0]_0 ));
  (* FSM_ENCODED_STATES = "WAIT_TMP:10,READ:11,IDLE:01,WAIT:00" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_fifo_state_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_0),
        .Q(fifo_state));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    broad_valid_i_1
       (.I0(broad_valid_i_2_n_0),
        .I1(broad_valid_i_3_n_0),
        .I2(broad_valid_i_4_n_0),
        .I3(broad_valid_i_5_n_0),
        .I4(broad_valid_i_6_n_0),
        .I5(broad_valid_i_7_n_0),
        .O(\da_addr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    broad_valid_i_10
       (.I0(da_addr[37]),
        .I1(da_addr[38]),
        .I2(da_addr[39]),
        .I3(da_addr[40]),
        .I4(da_addr[41]),
        .I5(da_addr[42]),
        .O(broad_valid_i_10_n_0));
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    broad_valid_i_2
       (.I0(broad_valid_i_8_n_0),
        .I1(da_addr[6]),
        .I2(da_addr[5]),
        .I3(da_addr[4]),
        .I4(broad_valid_i_9_n_0),
        .O(broad_valid_i_2_n_0));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    broad_valid_i_3
       (.I0(da_addr[22]),
        .I1(da_addr[23]),
        .I2(da_addr[24]),
        .I3(da_addr[21]),
        .I4(da_addr[19]),
        .I5(da_addr[20]),
        .O(broad_valid_i_3_n_0));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    broad_valid_i_4
       (.I0(da_addr[13]),
        .I1(da_addr[14]),
        .I2(da_addr[15]),
        .I3(da_addr[16]),
        .I4(da_addr[17]),
        .I5(da_addr[18]),
        .O(broad_valid_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    broad_valid_i_5
       (.I0(da_addr[47]),
        .I1(da_addr[46]),
        .I2(da_addr[45]),
        .I3(da_addr[44]),
        .I4(da_addr[43]),
        .I5(broad_valid_i_10_n_0),
        .O(broad_valid_i_5_n_0));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    broad_valid_i_6
       (.I0(da_addr[34]),
        .I1(da_addr[35]),
        .I2(da_addr[36]),
        .I3(da_addr[33]),
        .I4(da_addr[31]),
        .I5(da_addr[32]),
        .O(broad_valid_i_6_n_0));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    broad_valid_i_7
       (.I0(da_addr[25]),
        .I1(da_addr[26]),
        .I2(da_addr[27]),
        .I3(da_addr[28]),
        .I4(da_addr[29]),
        .I5(da_addr[30]),
        .O(broad_valid_i_7_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    broad_valid_i_8
       (.I0(da_addr[1]),
        .I1(da_addr[0]),
        .I2(da_addr[3]),
        .I3(da_addr[2]),
        .O(broad_valid_i_8_n_0));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    broad_valid_i_9
       (.I0(da_addr[10]),
        .I1(da_addr[11]),
        .I2(da_addr[12]),
        .I3(da_addr[9]),
        .I4(da_addr[7]),
        .I5(da_addr[8]),
        .O(broad_valid_i_9_n_0));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'h8B)) 
    \bytes_cnt[0]_i_1 
       (.I0(\terminator_location_reg[2]_0 [0]),
        .I1(get_terminator),
        .I2(\bytes_cnt_reg[1] [0]),
        .O(\terminator_location_reg[1]_0 [0]));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT4 #(
    .INIT(16'hB88B)) 
    \bytes_cnt[1]_i_1 
       (.I0(\terminator_location_reg[2]_0 [1]),
        .I1(get_terminator),
        .I2(\bytes_cnt_reg[1] [1]),
        .I3(\bytes_cnt_reg[1] [0]),
        .O(\terminator_location_reg[1]_0 [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \bytes_cnt[2]_i_1 
       (.I0(get_terminator),
        .I1(\bytes_cnt_reg[2] ),
        .O(get_terminator_reg_0));
  LUT2 #(
    .INIT(4'hB)) 
    check_reset_i_1
       (.I0(\FSM_sequential_fifo_state_reg[0]_0 ),
        .I1(fifo_state),
        .O(check_reset_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    check_reset_reg
       (.C(clk_i),
        .CE(check_reset_i_1_n_0),
        .CLR(reset_dcm),
        .D(check_reset_reg_0),
        .Q(check_reset));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[0] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[0]),
        .Q(da_addr[0]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[10] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[10]),
        .Q(da_addr[10]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[11] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[11]),
        .Q(da_addr[11]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[12] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[12]),
        .Q(da_addr[12]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[13] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[13]),
        .Q(da_addr[13]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[14] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[14]),
        .Q(da_addr[14]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[15] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[15]),
        .Q(da_addr[15]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[16] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[16]),
        .Q(da_addr[16]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[17] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[17]),
        .Q(da_addr[17]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[18] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[18]),
        .Q(da_addr[18]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[19] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[19]),
        .Q(da_addr[19]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[1] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[1]),
        .Q(da_addr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[20] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[20]),
        .Q(da_addr[20]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[21] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[21]),
        .Q(da_addr[21]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[22] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[22]),
        .Q(da_addr[22]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[23] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[23]),
        .Q(da_addr[23]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[24] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[24]),
        .Q(da_addr[24]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[25] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[25]),
        .Q(da_addr[25]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[26] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[26]),
        .Q(da_addr[26]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[27] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[27]),
        .Q(da_addr[27]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[28] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[28]),
        .Q(da_addr[28]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[29] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[29]),
        .Q(da_addr[29]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[2] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[2]),
        .Q(da_addr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[30] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[30]),
        .Q(da_addr[30]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[31] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[31]),
        .Q(da_addr[31]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[32] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[32]),
        .Q(da_addr[32]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[33] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[33]),
        .Q(da_addr[33]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[34] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[34]),
        .Q(da_addr[34]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[35] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[35]),
        .Q(da_addr[35]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[36] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[36]),
        .Q(da_addr[36]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[37] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[37]),
        .Q(da_addr[37]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[38] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[38]),
        .Q(da_addr[38]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[39] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[39]),
        .Q(da_addr[39]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[3] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[3]),
        .Q(da_addr[3]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[40] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[40]),
        .Q(da_addr[40]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[41] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[41]),
        .Q(da_addr[41]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[42] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[42]),
        .Q(da_addr[42]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[43] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[43]),
        .Q(da_addr[43]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[44] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[44]),
        .Q(da_addr[44]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[45] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[45]),
        .Q(da_addr[45]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[46] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[46]),
        .Q(da_addr[46]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[47] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[47]),
        .Q(da_addr[47]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[4] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[4]),
        .Q(da_addr[4]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[5] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[5]),
        .Q(da_addr[5]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[6] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[6]),
        .Q(da_addr[6]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[7] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[7]),
        .Q(da_addr[7]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[8] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[8]),
        .Q(da_addr[8]));
  FDCE #(
    .INIT(1'b0)) 
    \da_addr_reg[9] 
       (.C(clk_i),
        .CE(Q[0]),
        .CLR(reset_dcm),
        .D(rxd64_d1[9]),
        .Q(da_addr[9]));
  LUT6 #(
    .INIT(64'hFFFE000200020002)) 
    do_crc_check_i_1
       (.I0(get_terminator_d2),
        .I1(\terminator_location_reg[2]_0 [1]),
        .I2(\terminator_location_reg[2]_0 [0]),
        .I3(\terminator_location_reg[2]_0 [2]),
        .I4(wait_crc_check),
        .I5(do_crc_check_reg),
        .O(get_terminator_d2_reg));
  FDCE #(
    .INIT(1'b0)) 
    fifo_rd_en_reg
       (.C(clk_i),
        .CE(check_reset_i_1_n_0),
        .CLR(reset_dcm),
        .D(fifo_rd_en),
        .Q(fifo_rd_en_reg_n_0));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [0]),
        .Q(get_e_chk[0]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [1]),
        .Q(get_e_chk[1]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [2]),
        .Q(get_e_chk[2]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [3]),
        .Q(get_e_chk[3]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [4]),
        .Q(get_e_chk[4]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [5]),
        .Q(get_e_chk[5]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [6]),
        .Q(get_e_chk[6]));
  FDCE #(
    .INIT(1'b0)) 
    \get_e_chk_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\get_e_chk_reg[7]_0 [7]),
        .Q(get_e_chk[7]));
  LUT6 #(
    .INIT(64'h5555555555555554)) 
    get_error_code_i_1
       (.I0(get_error_code_reg_0),
        .I1(get_error_code_i_3_n_0),
        .I2(get_e_chk[4]),
        .I3(get_e_chk[6]),
        .I4(get_e_chk[1]),
        .I5(get_e_chk[3]),
        .O(get_error_code_i_1_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    get_error_code_i_3
       (.I0(get_e_chk[0]),
        .I1(get_e_chk[2]),
        .I2(get_e_chk[5]),
        .I3(get_e_chk[7]),
        .O(get_error_code_i_3_n_0));
  FDCE #(
    .INIT(1'b0)) 
    get_error_code_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(get_error_code_i_1_n_0),
        .Q(get_error_code));
  FDCE #(
    .INIT(1'b0)) 
    get_sfd_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(get_sfd0),
        .Q(get_sfd));
  FDCE #(
    .INIT(1'b0)) 
    get_terminator_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(E),
        .Q(get_terminator));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[0] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[40]),
        .Q(pad_remain0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[10] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[34]),
        .Q(\lt_data_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[11] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[35]),
        .Q(\lt_data_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[12] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[36]),
        .Q(\lt_data_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[13] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[37]),
        .Q(\lt_data_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[14] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[38]),
        .Q(\lt_data_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[15] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[39]),
        .Q(\lt_data_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[1] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[41]),
        .Q(\lt_data_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[2] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[42]),
        .Q(\lt_data_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[3] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[43]),
        .Q(\lt_data_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[4] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[44]),
        .Q(\lt_data_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[5] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[45]),
        .Q(\lt_data_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[6] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[46]),
        .Q(\lt_data_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[7] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[47]),
        .Q(\lt_data_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[8] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[32]),
        .Q(\lt_data_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \lt_data_reg[9] 
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(rxd64_d1[33]),
        .Q(\lt_data_reg_n_0_[9] ));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_1__0
       (.I0(rxc8_d3[0]),
        .I1(rxc_final[0]),
        .I2(inband_fcs),
        .O(vDataIn[0]));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_2
       (.I0(rxc8_d3[1]),
        .I1(rxc_final[1]),
        .I2(inband_fcs),
        .O(vDataIn[1]));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_3
       (.I0(rxc8_d3[2]),
        .I1(rxc_final[2]),
        .I2(inband_fcs),
        .O(vDataIn[2]));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_4
       (.I0(rxc8_d3[3]),
        .I1(rxc_final[3]),
        .I2(inband_fcs),
        .O(vDataIn[3]));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_5
       (.I0(rxc8_d3[4]),
        .I1(rxc_final[4]),
        .I2(inband_fcs),
        .O(vDataIn[4]));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_6
       (.I0(rxc8_d3[5]),
        .I1(rxc_final[5]),
        .I2(inband_fcs),
        .O(vDataIn[5]));
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_0_6_i_7
       (.I0(rxc8_d3[6]),
        .I1(rxc_final[6]),
        .I2(inband_fcs),
        .O(vDataIn[6]));
  LUT3 #(
    .INIT(8'h5C)) 
    mem_reg_0_63_7_7_i_1
       (.I0(rxc8_d3[7]),
        .I1(rxc_final[7]),
        .I2(inband_fcs),
        .O(vDataIn[7]));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    multi_valid_i_1
       (.I0(multi_valid_i_2_n_0),
        .I1(multi_valid_i_3_n_0),
        .I2(multi_valid_i_4_n_0),
        .I3(multi_valid_i_5_n_0),
        .I4(multi_valid_i_6_n_0),
        .I5(multi_valid_i_7_n_0),
        .O(\da_addr_reg[40]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    multi_valid_i_10
       (.I0(da_addr[37]),
        .I1(da_addr[35]),
        .I2(da_addr[36]),
        .I3(da_addr[42]),
        .I4(da_addr[38]),
        .I5(da_addr[41]),
        .O(multi_valid_i_10_n_0));
  LUT5 #(
    .INIT(32'hFFBFFFFF)) 
    multi_valid_i_2
       (.I0(multi_valid_i_8_n_0),
        .I1(da_addr[40]),
        .I2(da_addr[39]),
        .I3(da_addr[1]),
        .I4(multi_valid_i_9_n_0),
        .O(multi_valid_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    multi_valid_i_3
       (.I0(da_addr[19]),
        .I1(da_addr[17]),
        .I2(da_addr[18]),
        .I3(da_addr[14]),
        .I4(da_addr[15]),
        .I5(da_addr[16]),
        .O(multi_valid_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    multi_valid_i_4
       (.I0(da_addr[10]),
        .I1(da_addr[8]),
        .I2(da_addr[9]),
        .I3(da_addr[13]),
        .I4(da_addr[11]),
        .I5(da_addr[12]),
        .O(multi_valid_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    multi_valid_i_5
       (.I0(da_addr[45]),
        .I1(da_addr[44]),
        .I2(da_addr[43]),
        .I3(da_addr[47]),
        .I4(da_addr[46]),
        .I5(multi_valid_i_10_n_0),
        .O(multi_valid_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    multi_valid_i_6
       (.I0(da_addr[34]),
        .I1(da_addr[32]),
        .I2(da_addr[33]),
        .I3(da_addr[27]),
        .I4(da_addr[28]),
        .I5(da_addr[29]),
        .O(multi_valid_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    multi_valid_i_7
       (.I0(da_addr[22]),
        .I1(da_addr[20]),
        .I2(da_addr[21]),
        .I3(da_addr[26]),
        .I4(da_addr[23]),
        .I5(da_addr[24]),
        .O(multi_valid_i_7_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    multi_valid_i_8
       (.I0(da_addr[25]),
        .I1(da_addr[0]),
        .I2(da_addr[31]),
        .I3(da_addr[30]),
        .O(multi_valid_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    multi_valid_i_9
       (.I0(da_addr[7]),
        .I1(da_addr[5]),
        .I2(da_addr[6]),
        .I3(da_addr[2]),
        .I4(da_addr[3]),
        .I5(da_addr[4]),
        .O(multi_valid_i_9_n_0));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \pad_cnt[0]_i_1 
       (.I0(\pad_integer_reg_n_0_[0] ),
        .I1(\pad_cnt[2]_i_2_n_0 ),
        .O(pad_cnt[0]));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pad_cnt[1]_i_1 
       (.I0(\pad_cnt[2]_i_2_n_0 ),
        .I1(\pad_integer_reg_n_0_[1] ),
        .O(pad_cnt[1]));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT3 #(
    .INIT(8'h28)) 
    \pad_cnt[2]_i_1 
       (.I0(\pad_cnt[2]_i_2_n_0 ),
        .I1(\pad_integer_reg_n_0_[1] ),
        .I2(\pad_integer_reg_n_0_[2] ),
        .O(pad_cnt[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \pad_cnt[2]_i_2 
       (.I0(pad_remain0[0]),
        .I1(\lt_data_reg_n_0_[1] ),
        .I2(\lt_data_reg_n_0_[4] ),
        .I3(\lt_data_reg_n_0_[5] ),
        .I4(\lt_data_reg_n_0_[2] ),
        .I5(\lt_data_reg_n_0_[3] ),
        .O(\pad_cnt[2]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_cnt_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_cnt[0]),
        .Q(\pad_cnt_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_cnt_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_cnt[1]),
        .Q(\pad_cnt_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_cnt_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_cnt[2]),
        .Q(\pad_cnt_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_cnt_reg_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_3),
        .Q(pad_cnt_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_cnt_reg_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_2),
        .Q(pad_cnt_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_cnt_reg_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_1),
        .Q(pad_cnt_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    pad_frame_d1_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_6),
        .Q(pad_frame_d1_reg_n_0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    pad_frame_i_1
       (.I0(pad_frame_i_2_n_0),
        .I1(\lt_data_reg_n_0_[7] ),
        .I2(\lt_data_reg_n_0_[6] ),
        .I3(\lt_data_reg_n_0_[9] ),
        .I4(\lt_data_reg_n_0_[8] ),
        .I5(pad_frame_i_3_n_0),
        .O(pad_frame));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    pad_frame_i_2
       (.I0(\lt_data_reg_n_0_[12] ),
        .I1(\lt_data_reg_n_0_[13] ),
        .I2(\lt_data_reg_n_0_[10] ),
        .I3(\lt_data_reg_n_0_[11] ),
        .I4(\lt_data_reg_n_0_[15] ),
        .I5(\lt_data_reg_n_0_[14] ),
        .O(pad_frame_i_2_n_0));
  LUT6 #(
    .INIT(64'h33333FFF3333FFFE)) 
    pad_frame_i_3
       (.I0(pad_remain0[0]),
        .I1(\lt_data_reg_n_0_[5] ),
        .I2(\lt_data_reg_n_0_[2] ),
        .I3(\lt_data_reg_n_0_[3] ),
        .I4(\lt_data_reg_n_0_[4] ),
        .I5(\lt_data_reg_n_0_[1] ),
        .O(pad_frame_i_3_n_0));
  FDCE #(
    .INIT(1'b0)) 
    pad_frame_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_frame),
        .Q(pad_frame_reg_n_0));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'hC9)) 
    \pad_integer[0]_i_1 
       (.I0(\lt_data_reg_n_0_[2] ),
        .I1(\lt_data_reg_n_0_[3] ),
        .I2(\lt_data_reg_n_0_[1] ),
        .O(pad_integer1[3]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT4 #(
    .INIT(16'hCCC9)) 
    \pad_integer[1]_i_1 
       (.I0(\lt_data_reg_n_0_[1] ),
        .I1(\lt_data_reg_n_0_[4] ),
        .I2(\lt_data_reg_n_0_[2] ),
        .I3(\lt_data_reg_n_0_[3] ),
        .O(pad_integer1[4]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT5 #(
    .INIT(32'hAAAAAAA9)) 
    \pad_integer[2]_i_1 
       (.I0(\lt_data_reg_n_0_[5] ),
        .I1(\lt_data_reg_n_0_[2] ),
        .I2(\lt_data_reg_n_0_[3] ),
        .I3(\lt_data_reg_n_0_[4] ),
        .I4(\lt_data_reg_n_0_[1] ),
        .O(pad_integer1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_integer_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_integer1[3]),
        .Q(\pad_integer_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_integer_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_integer1[4]),
        .Q(\pad_integer_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_integer_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_integer1[5]),
        .Q(\pad_integer_reg_n_0_[2] ));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \pad_last_rxc[0]_i_1 
       (.I0(pad_remain[1]),
        .I1(pad_remain[0]),
        .I2(\pad_cnt[2]_i_2_n_0 ),
        .I3(pad_remain[2]),
        .O(pad_last_rxc[0]));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \pad_last_rxc[1]_i_1 
       (.I0(\pad_cnt[2]_i_2_n_0 ),
        .I1(pad_remain[2]),
        .I2(pad_remain[1]),
        .O(pad_last_rxc[1]));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT4 #(
    .INIT(16'hFF8F)) 
    \pad_last_rxc[2]_i_1 
       (.I0(pad_remain[1]),
        .I1(pad_remain[0]),
        .I2(\pad_cnt[2]_i_2_n_0 ),
        .I3(pad_remain[2]),
        .O(pad_last_rxc[2]));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \pad_last_rxc[3]_i_1 
       (.I0(pad_remain[2]),
        .I1(\pad_cnt[2]_i_2_n_0 ),
        .O(pad_last_rxc[3]));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT4 #(
    .INIT(16'hA8FF)) 
    \pad_last_rxc[4]_i_1 
       (.I0(pad_remain[2]),
        .I1(pad_remain[0]),
        .I2(pad_remain[1]),
        .I3(\pad_cnt[2]_i_2_n_0 ),
        .O(pad_last_rxc[4]));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'h8F)) 
    \pad_last_rxc[5]_i_1 
       (.I0(pad_remain[2]),
        .I1(pad_remain[1]),
        .I2(\pad_cnt[2]_i_2_n_0 ),
        .O(pad_last_rxc[5]));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT4 #(
    .INIT(16'h80FF)) 
    \pad_last_rxc[6]_i_1 
       (.I0(pad_remain[0]),
        .I1(pad_remain[1]),
        .I2(pad_remain[2]),
        .I3(\pad_cnt[2]_i_2_n_0 ),
        .O(pad_last_rxc[6]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[0]),
        .Q(\pad_last_rxc_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[1]),
        .Q(\pad_last_rxc_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[2]),
        .Q(\pad_last_rxc_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[3]),
        .Q(\pad_last_rxc_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[4]),
        .Q(\pad_last_rxc_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[5]),
        .Q(\pad_last_rxc_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \pad_last_rxc_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_last_rxc[6]),
        .Q(\pad_last_rxc_reg_n_0_[6] ));
  LUT1 #(
    .INIT(2'h1)) 
    \pad_remain[1]_i_1 
       (.I0(\lt_data_reg_n_0_[1] ),
        .O(pad_remain0[1]));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \pad_remain[2]_i_1 
       (.I0(\lt_data_reg_n_0_[1] ),
        .I1(\lt_data_reg_n_0_[2] ),
        .O(pad_remain0[2]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_remain_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_remain0[0]),
        .Q(pad_remain[0]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_remain_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_remain0[1]),
        .Q(pad_remain[1]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_remain_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(pad_remain0[2]),
        .Q(pad_remain[2]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[0] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[0] ),
        .Q(pad_rxc_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[1] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[1] ),
        .Q(pad_rxc_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[2] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[2] ),
        .Q(pad_rxc_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[3] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[3] ),
        .Q(pad_rxc_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[4] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[4] ),
        .Q(pad_rxc_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[5] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[5] ),
        .Q(pad_rxc_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \pad_rxc_reg_reg[6] 
       (.C(clk_i),
        .CE(pad_cnt_reg1),
        .CLR(reset_dcm),
        .D(\pad_last_rxc_reg_n_0_[6] ),
        .Q(pad_rxc_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    receiving_d1_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(receiving),
        .Q(in0));
  FDCE #(
    .INIT(1'b0)) 
    receiving_d2_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(in0),
        .Q(receiving_d2));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT3 #(
    .INIT(8'h02)) 
    rx_bad_frame_inferred_i_1
       (.I0(bad_frame_get),
        .I1(\FSM_sequential_fifo_state_reg[0]_0 ),
        .I2(fifo_state),
        .O(bad_frame_get_reg));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_70),
        .Q(\rx_data_reg[63]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_60),
        .Q(\rx_data_reg[63]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_59),
        .Q(\rx_data_reg[63]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_58),
        .Q(\rx_data_reg[63]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_57),
        .Q(\rx_data_reg[63]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_56),
        .Q(\rx_data_reg[63]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_55),
        .Q(\rx_data_reg[63]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_54),
        .Q(\rx_data_reg[63]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_53),
        .Q(\rx_data_reg[63]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_52),
        .Q(\rx_data_reg[63]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_51),
        .Q(\rx_data_reg[63]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_69),
        .Q(\rx_data_reg[63]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_50),
        .Q(\rx_data_reg[63]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_49),
        .Q(\rx_data_reg[63]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_48),
        .Q(\rx_data_reg[63]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_47),
        .Q(\rx_data_reg[63]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_46),
        .Q(\rx_data_reg[63]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_45),
        .Q(\rx_data_reg[63]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_44),
        .Q(\rx_data_reg[63]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_43),
        .Q(\rx_data_reg[63]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_42),
        .Q(\rx_data_reg[63]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_41),
        .Q(\rx_data_reg[63]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_68),
        .Q(\rx_data_reg[63]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_40),
        .Q(\rx_data_reg[63]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_39),
        .Q(\rx_data_reg[63]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_38),
        .Q(\rx_data_reg[63]_0 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_37),
        .Q(\rx_data_reg[63]_0 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_36),
        .Q(\rx_data_reg[63]_0 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_35),
        .Q(\rx_data_reg[63]_0 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_34),
        .Q(\rx_data_reg[63]_0 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_33),
        .Q(\rx_data_reg[63]_0 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_32),
        .Q(\rx_data_reg[63]_0 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_31),
        .Q(\rx_data_reg[63]_0 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_67),
        .Q(\rx_data_reg[63]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_30),
        .Q(\rx_data_reg[63]_0 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_29),
        .Q(\rx_data_reg[63]_0 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_28),
        .Q(\rx_data_reg[63]_0 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_27),
        .Q(\rx_data_reg[63]_0 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_26),
        .Q(\rx_data_reg[63]_0 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_25),
        .Q(\rx_data_reg[63]_0 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_24),
        .Q(\rx_data_reg[63]_0 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_23),
        .Q(\rx_data_reg[63]_0 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_22),
        .Q(\rx_data_reg[63]_0 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_21),
        .Q(\rx_data_reg[63]_0 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_66),
        .Q(\rx_data_reg[63]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_20),
        .Q(\rx_data_reg[63]_0 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_19),
        .Q(\rx_data_reg[63]_0 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_18),
        .Q(\rx_data_reg[63]_0 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_17),
        .Q(\rx_data_reg[63]_0 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_16),
        .Q(\rx_data_reg[63]_0 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_15),
        .Q(\rx_data_reg[63]_0 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_14),
        .Q(\rx_data_reg[63]_0 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_13),
        .Q(\rx_data_reg[63]_0 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_12),
        .Q(\rx_data_reg[63]_0 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_11),
        .Q(\rx_data_reg[63]_0 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_65),
        .Q(\rx_data_reg[63]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_10),
        .Q(\rx_data_reg[63]_0 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_9),
        .Q(\rx_data_reg[63]_0 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_8),
        .Q(\rx_data_reg[63]_0 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_7),
        .Q(\rx_data_reg[63]_0 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_64),
        .Q(\rx_data_reg[63]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_63),
        .Q(\rx_data_reg[63]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_62),
        .Q(\rx_data_reg[63]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxdatain_n_61),
        .Q(\rx_data_reg[63]_0 [9]));
  LUT2 #(
    .INIT(4'h1)) 
    \rx_data_valid[0]_i_2 
       (.I0(pad_cnt_reg[1]),
        .I1(pad_cnt_reg[2]),
        .O(\rx_data_valid[0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT4 #(
    .INIT(16'h10FF)) 
    \rx_data_valid[6]_i_2 
       (.I0(pad_cnt_reg[1]),
        .I1(pad_cnt_reg[2]),
        .I2(pad_frame_d1_reg_n_0),
        .I3(fifo_state),
        .O(\rx_data_valid[6]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    \rx_data_valid[6]_i_3 
       (.I0(pad_cnt_reg[2]),
        .I1(pad_cnt_reg[1]),
        .I2(pad_frame_d1_reg_n_0),
        .I3(fifo_state),
        .O(\rx_data_valid[6]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_10),
        .Q(\rx_data_valid_reg[7]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_9),
        .Q(\rx_data_valid_reg[7]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_8),
        .Q(\rx_data_valid_reg[7]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_7),
        .Q(\rx_data_valid_reg[7]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_6),
        .Q(\rx_data_valid_reg[7]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_5),
        .Q(\rx_data_valid_reg[7]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_4),
        .Q(\rx_data_valid_reg[7]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \rx_data_valid_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxcntrlin_n_3),
        .Q(\rx_data_valid_reg[7]_0 [7]));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT3 #(
    .INIT(8'h02)) 
    rx_good_frame_inferred_i_1
       (.I0(good_frame_get),
        .I1(\FSM_sequential_fifo_state_reg[0]_0 ),
        .I2(fifo_state),
        .O(good_frame_get_reg));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[64]),
        .Q(rxc8_d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[65]),
        .Q(rxc8_d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[66]),
        .Q(rxc8_d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[67]),
        .Q(rxc8_d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[68]),
        .Q(rxc8_d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[69]),
        .Q(rxc8_d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[70]),
        .Q(rxc8_d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[71]),
        .Q(rxc8_d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[0]),
        .Q(rxc8_d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[1]),
        .Q(rxc8_d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[2]),
        .Q(rxc8_d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[3]),
        .Q(rxc8_d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[4]),
        .Q(rxc8_d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[5]),
        .Q(rxc8_d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[6]),
        .Q(rxc8_d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d1[7]),
        .Q(rxc8_d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[0]),
        .Q(rxc8_d3[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[1]),
        .Q(rxc8_d3[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[2]),
        .Q(rxc8_d3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[3]),
        .Q(rxc8_d3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[4]),
        .Q(rxc8_d3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[5]),
        .Q(rxc8_d3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[6]),
        .Q(rxc8_d3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_d3_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxc8_d2[7]),
        .Q(rxc8_d3[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(1'b1),
        .Q(rxc_end_data[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(D[0]),
        .Q(rxc_end_data[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(D[1]),
        .Q(rxc_end_data[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[4] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(D[2]),
        .Q(rxc_end_data[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[5] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(D[3]),
        .Q(rxc_end_data[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[6] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(D[4]),
        .Q(rxc_end_data[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_end_data_reg[7] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(D[5]),
        .Q(rxc_end_data[7]));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[0]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[0]),
        .O(\rxc_final[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[1]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[1]),
        .O(\rxc_final[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[2]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[2]),
        .O(\rxc_final[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hF100F111)) 
    \rxc_final[3]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .O(\rxc_final[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[4]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[4]),
        .O(\rxc_final[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[5]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[5]),
        .O(\rxc_final[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[6]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[6]),
        .O(\rxc_final[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFF11101000111)) 
    \rxc_final[7]_i_1 
       (.I0(get_error_code),
        .I1(get_error_code_reg_0),
        .I2(get_terminator),
        .I3(this_cycle_reg_n_0),
        .I4(get_terminator_d1),
        .I5(rxc_end_data[7]),
        .O(\rxc_final[7]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[0]_i_1_n_0 ),
        .Q(rxc_final[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[1]_i_1_n_0 ),
        .Q(rxc_final[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[2]_i_1_n_0 ),
        .Q(rxc_final[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[3]_i_1_n_0 ),
        .Q(rxc_final[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[4]_i_1_n_0 ),
        .Q(rxc_final[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[5]_i_1_n_0 ),
        .Q(rxc_final[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[6]_i_1_n_0 ),
        .Q(rxc_final[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc_final_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\rxc_final[7]_i_1_n_0 ),
        .Q(rxc_final[7]));
  switch_elements_SwitchSyncFIFO__parameterized0 rxcntrlin
       (.D({rxcntrlin_n_0,rxcntrlin_n_1}),
        .Q({fifo_state,\FSM_sequential_fifo_state_reg[0]_0 }),
        .bad_frame_get(bad_frame_get),
        .clk_i(clk_i),
        .good_frame_get(good_frame_get),
        .\ovDataOut_reg[5]_0 (rxcntrlin_n_2),
        .\ovDataOut_reg[7]_0 ({rxcntrlin_n_3,rxcntrlin_n_4,rxcntrlin_n_5,rxcntrlin_n_6,rxcntrlin_n_7,rxcntrlin_n_8,rxcntrlin_n_9,rxcntrlin_n_10}),
        .\qvRAddr_reg[6] (fifo_rd_en_reg_n_0),
        .receiving_d2(receiving_d2),
        .reset_dcm(reset_dcm),
        .\rx_data_valid_reg[0] (\rx_data_valid[0]_i_2_n_0 ),
        .\rx_data_valid_reg[1] (\rx_data_valid[6]_i_2_n_0 ),
        .\rx_data_valid_reg[1]_0 (\rx_data_valid[6]_i_3_n_0 ),
        .\rx_data_valid_reg[6] (pad_rxc_reg),
        .\rx_data_valid_reg[7] (pad_cnt_reg),
        .\rx_data_valid_reg[7]_0 (pad_frame_d1_reg_n_0),
        .rxfifo_empty(rxfifo_empty),
        .vDataIn(vDataIn));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[0]),
        .Q(rxd64_d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[10]),
        .Q(rxd64_d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[11]),
        .Q(rxd64_d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[12]),
        .Q(rxd64_d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[13]),
        .Q(rxd64_d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[14]),
        .Q(rxd64_d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[15]),
        .Q(rxd64_d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[16]),
        .Q(rxd64_d1[16]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[17]),
        .Q(rxd64_d1[17]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[18]),
        .Q(rxd64_d1[18]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[19]),
        .Q(rxd64_d1[19]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[1]),
        .Q(rxd64_d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[20]),
        .Q(rxd64_d1[20]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[21]),
        .Q(rxd64_d1[21]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[22]),
        .Q(rxd64_d1[22]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[23]),
        .Q(rxd64_d1[23]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[24]),
        .Q(rxd64_d1[24]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[25]),
        .Q(rxd64_d1[25]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[26]),
        .Q(rxd64_d1[26]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[27]),
        .Q(rxd64_d1[27]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[28]),
        .Q(rxd64_d1[28]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[29]),
        .Q(rxd64_d1[29]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[2]),
        .Q(rxd64_d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[30]),
        .Q(rxd64_d1[30]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[31]),
        .Q(rxd64_d1[31]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[32]),
        .Q(rxd64_d1[32]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[33]),
        .Q(rxd64_d1[33]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[34]),
        .Q(rxd64_d1[34]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[35]),
        .Q(rxd64_d1[35]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[36]),
        .Q(rxd64_d1[36]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[37]),
        .Q(rxd64_d1[37]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[38]),
        .Q(rxd64_d1[38]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[39]),
        .Q(rxd64_d1[39]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[3]),
        .Q(rxd64_d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[40]),
        .Q(rxd64_d1[40]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[41]),
        .Q(rxd64_d1[41]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[42]),
        .Q(rxd64_d1[42]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[43]),
        .Q(rxd64_d1[43]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[44]),
        .Q(rxd64_d1[44]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[45]),
        .Q(rxd64_d1[45]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[46]),
        .Q(rxd64_d1[46]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[47]),
        .Q(rxd64_d1[47]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[48]),
        .Q(rxd64_d1[48]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[49]),
        .Q(rxd64_d1[49]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[4]),
        .Q(rxd64_d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[50]),
        .Q(rxd64_d1[50]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[51]),
        .Q(rxd64_d1[51]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[52]),
        .Q(rxd64_d1[52]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[53]),
        .Q(rxd64_d1[53]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[54]),
        .Q(rxd64_d1[54]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[55]),
        .Q(rxd64_d1[55]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[56]),
        .Q(rxd64_d1[56]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[57]),
        .Q(rxd64_d1[57]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[58]),
        .Q(rxd64_d1[58]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[59]),
        .Q(rxd64_d1[59]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[5]),
        .Q(rxd64_d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[60]),
        .Q(rxd64_d1[60]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[61]),
        .Q(rxd64_d1[61]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[62]),
        .Q(rxd64_d1[62]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[63]),
        .Q(rxd64_d1[63]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[6]),
        .Q(rxd64_d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[7]),
        .Q(rxd64_d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[8]),
        .Q(rxd64_d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(qvDataOut[9]),
        .Q(rxd64_d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[0]),
        .Q(rxd64_d2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[10]),
        .Q(rxd64_d2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[11]),
        .Q(rxd64_d2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[12]),
        .Q(rxd64_d2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[13]),
        .Q(rxd64_d2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[14]),
        .Q(rxd64_d2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[15]),
        .Q(rxd64_d2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[16]),
        .Q(rxd64_d2[16]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[17]),
        .Q(rxd64_d2[17]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[18]),
        .Q(rxd64_d2[18]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[19]),
        .Q(rxd64_d2[19]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[1]),
        .Q(rxd64_d2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[20]),
        .Q(rxd64_d2[20]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[21]),
        .Q(rxd64_d2[21]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[22]),
        .Q(rxd64_d2[22]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[23]),
        .Q(rxd64_d2[23]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[24]),
        .Q(rxd64_d2[24]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[25]),
        .Q(rxd64_d2[25]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[26]),
        .Q(rxd64_d2[26]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[27]),
        .Q(rxd64_d2[27]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[28]),
        .Q(rxd64_d2[28]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[29]),
        .Q(rxd64_d2[29]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[2]),
        .Q(rxd64_d2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[30]),
        .Q(rxd64_d2[30]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[31]),
        .Q(rxd64_d2[31]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[32]),
        .Q(rxd64_d2[32]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[33]),
        .Q(rxd64_d2[33]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[34]),
        .Q(rxd64_d2[34]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[35]),
        .Q(rxd64_d2[35]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[36]),
        .Q(rxd64_d2[36]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[37]),
        .Q(rxd64_d2[37]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[38]),
        .Q(rxd64_d2[38]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[39]),
        .Q(rxd64_d2[39]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[3]),
        .Q(rxd64_d2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[40]),
        .Q(rxd64_d2[40]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[41]),
        .Q(rxd64_d2[41]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[42]),
        .Q(rxd64_d2[42]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[43]),
        .Q(rxd64_d2[43]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[44]),
        .Q(rxd64_d2[44]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[45]),
        .Q(rxd64_d2[45]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[46]),
        .Q(rxd64_d2[46]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[47]),
        .Q(rxd64_d2[47]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[48]),
        .Q(rxd64_d2[48]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[49]),
        .Q(rxd64_d2[49]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[4]),
        .Q(rxd64_d2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[50]),
        .Q(rxd64_d2[50]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[51]),
        .Q(rxd64_d2[51]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[52]),
        .Q(rxd64_d2[52]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[53]),
        .Q(rxd64_d2[53]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[54]),
        .Q(rxd64_d2[54]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[55]),
        .Q(rxd64_d2[55]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[56]),
        .Q(rxd64_d2[56]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[57]),
        .Q(rxd64_d2[57]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[58]),
        .Q(rxd64_d2[58]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[59]),
        .Q(rxd64_d2[59]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[5]),
        .Q(rxd64_d2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[60]),
        .Q(rxd64_d2[60]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[61]),
        .Q(rxd64_d2[61]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[62]),
        .Q(rxd64_d2[62]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[63]),
        .Q(rxd64_d2[63]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[6]),
        .Q(rxd64_d2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[7]),
        .Q(rxd64_d2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[8]),
        .Q(rxd64_d2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d1[9]),
        .Q(rxd64_d2[9]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[0]),
        .Q(rxd64_d3[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[10]),
        .Q(rxd64_d3[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[11]),
        .Q(rxd64_d3[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[12]),
        .Q(rxd64_d3[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[13]),
        .Q(rxd64_d3[13]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[14]),
        .Q(rxd64_d3[14]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[15]),
        .Q(rxd64_d3[15]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[16]),
        .Q(rxd64_d3[16]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[17]),
        .Q(rxd64_d3[17]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[18]),
        .Q(rxd64_d3[18]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[19]),
        .Q(rxd64_d3[19]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[1]),
        .Q(rxd64_d3[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[20]),
        .Q(rxd64_d3[20]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[21]),
        .Q(rxd64_d3[21]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[22]),
        .Q(rxd64_d3[22]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[23]),
        .Q(rxd64_d3[23]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[24]),
        .Q(rxd64_d3[24]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[25]),
        .Q(rxd64_d3[25]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[26]),
        .Q(rxd64_d3[26]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[27]),
        .Q(rxd64_d3[27]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[28]),
        .Q(rxd64_d3[28]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[29]),
        .Q(rxd64_d3[29]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[2]),
        .Q(rxd64_d3[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[30]),
        .Q(rxd64_d3[30]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[31]),
        .Q(rxd64_d3[31]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[32]),
        .Q(rxd64_d3[32]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[33]),
        .Q(rxd64_d3[33]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[34]),
        .Q(rxd64_d3[34]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[35]),
        .Q(rxd64_d3[35]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[36]),
        .Q(rxd64_d3[36]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[37]),
        .Q(rxd64_d3[37]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[38]),
        .Q(rxd64_d3[38]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[39]),
        .Q(rxd64_d3[39]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[3]),
        .Q(rxd64_d3[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[40]),
        .Q(rxd64_d3[40]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[41]),
        .Q(rxd64_d3[41]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[42]),
        .Q(rxd64_d3[42]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[43]),
        .Q(rxd64_d3[43]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[44]),
        .Q(rxd64_d3[44]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[45]),
        .Q(rxd64_d3[45]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[46]),
        .Q(rxd64_d3[46]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[47]),
        .Q(rxd64_d3[47]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[48]),
        .Q(rxd64_d3[48]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[49]),
        .Q(rxd64_d3[49]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[4]),
        .Q(rxd64_d3[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[50]),
        .Q(rxd64_d3[50]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[51]),
        .Q(rxd64_d3[51]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[52]),
        .Q(rxd64_d3[52]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[53]),
        .Q(rxd64_d3[53]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[54]),
        .Q(rxd64_d3[54]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[55]),
        .Q(rxd64_d3[55]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[56]),
        .Q(rxd64_d3[56]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[57]),
        .Q(rxd64_d3[57]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[58]),
        .Q(rxd64_d3[58]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[59]),
        .Q(rxd64_d3[59]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[5]),
        .Q(rxd64_d3[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[60]),
        .Q(rxd64_d3[60]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[61]),
        .Q(rxd64_d3[61]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[62]),
        .Q(rxd64_d3[62]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[63]),
        .Q(rxd64_d3[63]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[6]),
        .Q(rxd64_d3[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[7]),
        .Q(rxd64_d3[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[8]),
        .Q(rxd64_d3[8]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_d3_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(rxd64_d2[9]),
        .Q(rxd64_d3[9]));
  switch_elements_SwitchSyncFIFO rxdatain
       (.D({rxdatain_n_1,rxdatain_n_2,rxdatain_n_3}),
        .Q({\pad_cnt_reg_n_0_[2] ,\pad_cnt_reg_n_0_[1] ,\pad_cnt_reg_n_0_[0] }),
        .clk_i(clk_i),
        .fifo_rd_en(fifo_rd_en),
        .fifo_rd_en_reg({fifo_state,\FSM_sequential_fifo_state_reg[0]_0 }),
        .fifo_rd_en_reg_0(rxcntrlin_n_2),
        .\ovDataOut_reg[63]_0 ({rxdatain_n_7,rxdatain_n_8,rxdatain_n_9,rxdatain_n_10,rxdatain_n_11,rxdatain_n_12,rxdatain_n_13,rxdatain_n_14,rxdatain_n_15,rxdatain_n_16,rxdatain_n_17,rxdatain_n_18,rxdatain_n_19,rxdatain_n_20,rxdatain_n_21,rxdatain_n_22,rxdatain_n_23,rxdatain_n_24,rxdatain_n_25,rxdatain_n_26,rxdatain_n_27,rxdatain_n_28,rxdatain_n_29,rxdatain_n_30,rxdatain_n_31,rxdatain_n_32,rxdatain_n_33,rxdatain_n_34,rxdatain_n_35,rxdatain_n_36,rxdatain_n_37,rxdatain_n_38,rxdatain_n_39,rxdatain_n_40,rxdatain_n_41,rxdatain_n_42,rxdatain_n_43,rxdatain_n_44,rxdatain_n_45,rxdatain_n_46,rxdatain_n_47,rxdatain_n_48,rxdatain_n_49,rxdatain_n_50,rxdatain_n_51,rxdatain_n_52,rxdatain_n_53,rxdatain_n_54,rxdatain_n_55,rxdatain_n_56,rxdatain_n_57,rxdatain_n_58,rxdatain_n_59,rxdatain_n_60,rxdatain_n_61,rxdatain_n_62,rxdatain_n_63,rxdatain_n_64,rxdatain_n_65,rxdatain_n_66,rxdatain_n_67,rxdatain_n_68,rxdatain_n_69,rxdatain_n_70}),
        .pad_cnt_reg1(pad_cnt_reg1),
        .\pad_cnt_reg_reg[0] (pad_cnt_reg),
        .pad_frame_d1_reg(pad_frame_d1_reg_n_0),
        .\pad_rxc_reg_reg[0] (pad_frame_reg_n_0),
        .qEmpty_reg(rxdatain_n_6),
        .\qvRAddr_reg[6] (fifo_rd_en_reg_n_0),
        .receiving_d2(receiving_d2),
        .reset_dcm(reset_dcm),
        .rxd64_d3(rxd64_d3),
        .rxfifo_empty(rxfifo_empty));
  FDCE #(
    .INIT(1'b0)) 
    tagged_frame_reg
       (.C(clk_i),
        .CE(Q[1]),
        .CLR(reset_dcm),
        .D(tagged_frame_reg_0),
        .Q(tagged_frame));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_location_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(\terminator_location_reg[2]_1 [0]),
        .Q(\terminator_location_reg[2]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_location_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(\terminator_location_reg[2]_1 [1]),
        .Q(\terminator_location_reg[2]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \terminator_location_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(\terminator_location_reg[2]_1 [2]),
        .Q(\terminator_location_reg[2]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    this_cycle_reg
       (.C(clk_i),
        .CE(E),
        .CLR(reset_dcm),
        .D(this_cycle),
        .Q(this_cycle_reg_n_0));
endmodule

(* ORIG_REF_NAME = "rxLenTypChecker" *) 
module switch_elements_rxLenTypChecker
   (large_error,
    small_error,
    padded_frame,
    length_65_127,
    length_128_255,
    length_256_511,
    length_512_1023,
    jumbo_frame,
    D,
    bad_frame_get0,
    \location_reg_reg[0]_0 ,
    \location_reg_reg[2]_0 ,
    \location_reg_reg[0]_1 ,
    large_error_reg_0,
    clk_i,
    reset_dcm,
    small_error0,
    padded_frame0,
    length_65_1270,
    length_128_2550,
    length_256_5110,
    length_512_10230,
    jumbo_frame0,
    get_error_code,
    Q,
    get_terminator,
    bad_frame_get_reg,
    vlan_enable,
    tagged_frame,
    large_error_i_4,
    large_error_i_4_0,
    jumbo_enable,
    large_error_reg_1,
    large_error_reg_2,
    \location_reg_reg[2]_1 );
  output large_error;
  output small_error;
  output padded_frame;
  output length_65_127;
  output length_128_255;
  output length_256_511;
  output length_512_1023;
  output jumbo_frame;
  output [1:0]D;
  output bad_frame_get0;
  output \location_reg_reg[0]_0 ;
  output [0:0]\location_reg_reg[2]_0 ;
  output \location_reg_reg[0]_1 ;
  input large_error_reg_0;
  input clk_i;
  input reset_dcm;
  input small_error0;
  input padded_frame0;
  input length_65_1270;
  input length_128_2550;
  input length_256_5110;
  input length_512_10230;
  input jumbo_frame0;
  input get_error_code;
  input [1:0]Q;
  input get_terminator;
  input [0:0]bad_frame_get_reg;
  input vlan_enable;
  input tagged_frame;
  input large_error_i_4;
  input large_error_i_4_0;
  input jumbo_enable;
  input large_error_reg_1;
  input large_error_reg_2;
  input [2:0]\location_reg_reg[2]_1 ;

  wire [1:0]D;
  wire [1:0]Q;
  wire bad_frame_get0;
  wire [0:0]bad_frame_get_reg;
  wire clk_i;
  wire get_error_code;
  wire get_terminator;
  wire jumbo_enable;
  wire jumbo_frame;
  wire jumbo_frame0;
  wire large_error;
  wire large_error_i_4;
  wire large_error_i_4_0;
  wire large_error_reg_0;
  wire large_error_reg_1;
  wire large_error_reg_2;
  wire length_128_255;
  wire length_128_2550;
  wire length_256_511;
  wire length_256_5110;
  wire length_512_1023;
  wire length_512_10230;
  wire length_65_127;
  wire length_65_1270;
  wire [1:0]location_reg;
  wire \location_reg_reg[0]_0 ;
  wire \location_reg_reg[0]_1 ;
  wire [0:0]\location_reg_reg[2]_0 ;
  wire [2:0]\location_reg_reg[2]_1 ;
  wire padded_frame;
  wire padded_frame0;
  wire reset_dcm;
  wire small_error;
  wire small_error0;
  wire tagged_frame;
  wire vlan_enable;

  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT4 #(
    .INIT(16'hAAA8)) 
    \FSM_onehot_rxstate_next_reg[4]_i_1 
       (.I0(Q[0]),
        .I1(large_error),
        .I2(small_error),
        .I3(get_error_code),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT5 #(
    .INIT(32'h01000000)) 
    \FSM_onehot_rxstate_next_reg[5]_i_1 
       (.I0(large_error),
        .I1(small_error),
        .I2(get_error_code),
        .I3(Q[0]),
        .I4(get_terminator),
        .O(D[1]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    bad_frame_get_i_1
       (.I0(Q[1]),
        .I1(large_error),
        .I2(small_error),
        .I3(bad_frame_get_reg),
        .O(bad_frame_get0));
  FDCE #(
    .INIT(1'b0)) 
    jumbo_frame_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(jumbo_frame0),
        .Q(jumbo_frame));
  LUT6 #(
    .INIT(64'hFF00FF00FF000707)) 
    large_error_i_2
       (.I0(location_reg[0]),
        .I1(location_reg[1]),
        .I2(\location_reg_reg[2]_0 ),
        .I3(jumbo_enable),
        .I4(large_error_reg_1),
        .I5(large_error_reg_2),
        .O(\location_reg_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF777)) 
    large_error_i_8
       (.I0(location_reg[0]),
        .I1(location_reg[1]),
        .I2(vlan_enable),
        .I3(tagged_frame),
        .I4(large_error_i_4),
        .I5(large_error_i_4_0),
        .O(\location_reg_reg[0]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    large_error_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(large_error_reg_0),
        .Q(large_error));
  FDCE #(
    .INIT(1'b0)) 
    length_128_255_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(length_128_2550),
        .Q(length_128_255));
  FDCE #(
    .INIT(1'b0)) 
    length_256_511_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(length_256_5110),
        .Q(length_256_511));
  FDCE #(
    .INIT(1'b0)) 
    length_512_1023_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(length_512_10230),
        .Q(length_512_1023));
  FDCE #(
    .INIT(1'b0)) 
    length_65_127_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(length_65_1270),
        .Q(length_65_127));
  FDCE #(
    .INIT(1'b0)) 
    \location_reg_reg[0] 
       (.C(clk_i),
        .CE(get_terminator),
        .CLR(reset_dcm),
        .D(\location_reg_reg[2]_1 [0]),
        .Q(location_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \location_reg_reg[1] 
       (.C(clk_i),
        .CE(get_terminator),
        .CLR(reset_dcm),
        .D(\location_reg_reg[2]_1 [1]),
        .Q(location_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \location_reg_reg[2] 
       (.C(clk_i),
        .CE(get_terminator),
        .CLR(reset_dcm),
        .D(\location_reg_reg[2]_1 [2]),
        .Q(\location_reg_reg[2]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    padded_frame_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(padded_frame0),
        .Q(padded_frame));
  FDCE #(
    .INIT(1'b0)) 
    small_error_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(small_error0),
        .Q(small_error));
endmodule

(* ORIG_REF_NAME = "rxLinkFaultState" *) 
module switch_elements_rxLinkFaultState
   (Q,
    \link_fault_reg[1]_0 ,
    remote_fault,
    rxclk_180,
    AR,
    \FSM_sequential_linkstate_reg[0]_0 ,
    local_fault);
  output [0:0]Q;
  output [1:0]\link_fault_reg[1]_0 ;
  input remote_fault;
  input rxclk_180;
  input [0:0]AR;
  input \FSM_sequential_linkstate_reg[0]_0 ;
  input local_fault;

  wire [0:0]AR;
  wire \FSM_sequential_linkstate[0]_i_1_n_0 ;
  wire \FSM_sequential_linkstate[0]_i_2_n_0 ;
  wire \FSM_sequential_linkstate[0]_i_3_n_0 ;
  wire \FSM_sequential_linkstate[1]_i_1_n_0 ;
  wire \FSM_sequential_linkstate[1]_i_2_n_0 ;
  wire \FSM_sequential_linkstate_reg[0]_0 ;
  wire [0:0]Q;
  wire \col_cnt[2]_i_1_n_0 ;
  wire \col_cnt[3]_i_1_n_0 ;
  wire \col_cnt[4]_i_1_n_0 ;
  wire [5:0]col_cnt_reg;
  wire [0:0]last_seq_type;
  wire [0:0]link_fault0_in;
  wire \link_fault[1]_i_1_n_0 ;
  wire [1:0]\link_fault_reg[1]_0 ;
  wire [0:0]linkstate;
  wire local_fault;
  wire [5:0]p_0_in__6;
  wire remote_fault;
  wire reset_col_cnt;
  wire reset_col_cnt_0;
  wire rxclk_180;
  wire seq_cnt_i_1_n_0;
  wire seq_cnt_reg_n_0;
  wire [0:0]seq_type;

  LUT6 #(
    .INIT(64'h000F777FFFFF0000)) 
    \FSM_sequential_linkstate[0]_i_1 
       (.I0(\FSM_sequential_linkstate[0]_i_2_n_0 ),
        .I1(col_cnt_reg[5]),
        .I2(\FSM_sequential_linkstate[0]_i_3_n_0 ),
        .I3(seq_cnt_reg_n_0),
        .I4(\FSM_sequential_linkstate_reg[0]_0 ),
        .I5(linkstate),
        .O(\FSM_sequential_linkstate[0]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \FSM_sequential_linkstate[0]_i_2 
       (.I0(col_cnt_reg[4]),
        .I1(col_cnt_reg[3]),
        .I2(col_cnt_reg[1]),
        .I3(col_cnt_reg[0]),
        .I4(col_cnt_reg[2]),
        .O(\FSM_sequential_linkstate[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF666F)) 
    \FSM_sequential_linkstate[0]_i_3 
       (.I0(last_seq_type),
        .I1(seq_type),
        .I2(remote_fault),
        .I3(local_fault),
        .I4(Q),
        .O(\FSM_sequential_linkstate[0]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \FSM_sequential_linkstate[1]_i_1 
       (.I0(Q),
        .I1(linkstate),
        .O(\FSM_sequential_linkstate[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0060006000600000)) 
    \FSM_sequential_linkstate[1]_i_2 
       (.I0(last_seq_type),
        .I1(seq_type),
        .I2(linkstate),
        .I3(Q),
        .I4(local_fault),
        .I5(remote_fault),
        .O(\FSM_sequential_linkstate[1]_i_2_n_0 ));
  (* FSM_ENCODED_STATES = "IDLE:00,LinkFaultDetect:01,NewFaultType:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_linkstate_reg[0] 
       (.C(rxclk_180),
        .CE(\FSM_sequential_linkstate[1]_i_1_n_0 ),
        .CLR(AR),
        .D(\FSM_sequential_linkstate[0]_i_1_n_0 ),
        .Q(linkstate));
  (* FSM_ENCODED_STATES = "IDLE:00,LinkFaultDetect:01,NewFaultType:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_linkstate_reg[1] 
       (.C(rxclk_180),
        .CE(\FSM_sequential_linkstate[1]_i_1_n_0 ),
        .CLR(AR),
        .D(\FSM_sequential_linkstate[1]_i_2_n_0 ),
        .Q(Q));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \col_cnt[0]_i_1 
       (.I0(col_cnt_reg[0]),
        .I1(reset_col_cnt),
        .O(p_0_in__6[0]));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \col_cnt[1]_i_1 
       (.I0(col_cnt_reg[1]),
        .I1(col_cnt_reg[0]),
        .I2(reset_col_cnt),
        .O(p_0_in__6[1]));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT4 #(
    .INIT(16'h1540)) 
    \col_cnt[2]_i_1 
       (.I0(reset_col_cnt),
        .I1(col_cnt_reg[0]),
        .I2(col_cnt_reg[1]),
        .I3(col_cnt_reg[2]),
        .O(\col_cnt[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT5 #(
    .INIT(32'h15554000)) 
    \col_cnt[3]_i_1 
       (.I0(reset_col_cnt),
        .I1(col_cnt_reg[1]),
        .I2(col_cnt_reg[0]),
        .I3(col_cnt_reg[2]),
        .I4(col_cnt_reg[3]),
        .O(\col_cnt[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    \col_cnt[4]_i_1 
       (.I0(reset_col_cnt),
        .I1(col_cnt_reg[2]),
        .I2(col_cnt_reg[0]),
        .I3(col_cnt_reg[1]),
        .I4(col_cnt_reg[3]),
        .I5(col_cnt_reg[4]),
        .O(\col_cnt[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \col_cnt[5]_i_1 
       (.I0(\FSM_sequential_linkstate[0]_i_2_n_0 ),
        .I1(col_cnt_reg[5]),
        .I2(reset_col_cnt),
        .O(p_0_in__6[5]));
  FDCE #(
    .INIT(1'b0)) 
    \col_cnt_reg[0] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(p_0_in__6[0]),
        .Q(col_cnt_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \col_cnt_reg[1] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(p_0_in__6[1]),
        .Q(col_cnt_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \col_cnt_reg[2] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(\col_cnt[2]_i_1_n_0 ),
        .Q(col_cnt_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \col_cnt_reg[3] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(\col_cnt[3]_i_1_n_0 ),
        .Q(col_cnt_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \col_cnt_reg[4] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(\col_cnt[4]_i_1_n_0 ),
        .Q(col_cnt_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \col_cnt_reg[5] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(p_0_in__6[5]),
        .Q(col_cnt_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \last_seq_type_reg[0] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(seq_type),
        .Q(last_seq_type));
  LUT3 #(
    .INIT(8'h08)) 
    \link_fault[0]_i_1 
       (.I0(seq_type),
        .I1(linkstate),
        .I2(Q),
        .O(link_fault0_in));
  LUT4 #(
    .INIT(16'h1F11)) 
    \link_fault[1]_i_1 
       (.I0(linkstate),
        .I1(Q),
        .I2(\FSM_sequential_linkstate[0]_i_3_n_0 ),
        .I3(seq_cnt_reg_n_0),
        .O(\link_fault[1]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \link_fault_reg[0] 
       (.C(rxclk_180),
        .CE(\link_fault[1]_i_1_n_0 ),
        .CLR(AR),
        .D(link_fault0_in),
        .Q(\link_fault_reg[1]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \link_fault_reg[1] 
       (.C(rxclk_180),
        .CE(\link_fault[1]_i_1_n_0 ),
        .CLR(AR),
        .D(1'b0),
        .Q(\link_fault_reg[1]_0 [1]));
  LUT4 #(
    .INIT(16'h55FD)) 
    reset_col_cnt_i_1
       (.I0(linkstate),
        .I1(remote_fault),
        .I2(local_fault),
        .I3(Q),
        .O(reset_col_cnt_0));
  FDPE #(
    .INIT(1'b1)) 
    reset_col_cnt_reg
       (.C(rxclk_180),
        .CE(\FSM_sequential_linkstate[1]_i_1_n_0 ),
        .D(reset_col_cnt_0),
        .PRE(AR),
        .Q(reset_col_cnt));
  LUT3 #(
    .INIT(8'hD0)) 
    seq_cnt_i_1
       (.I0(\FSM_sequential_linkstate[0]_i_3_n_0 ),
        .I1(seq_cnt_reg_n_0),
        .I2(linkstate),
        .O(seq_cnt_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    seq_cnt_reg
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(seq_cnt_i_1_n_0),
        .Q(seq_cnt_reg_n_0));
  FDCE #(
    .INIT(1'b0)) 
    \seq_type_reg[0] 
       (.C(rxclk_180),
        .CE(1'b1),
        .CLR(AR),
        .D(remote_fault),
        .Q(seq_type));
endmodule

(* ORIG_REF_NAME = "rxNumCounter" *) 
module switch_elements_rxNumCounter
   (\value_reg[10] ,
    \value_reg[9] ,
    \value_reg[11] ,
    \value_reg[2] ,
    jumbo_frame0,
    \value_reg[8] ,
    \value_reg[4] ,
    \value_reg[1] ,
    \value_reg[1]_0 ,
    length_256_5110,
    length_512_10230,
    length_65_1270,
    padded_frame0,
    small_error0,
    length_128_2550,
    \value_reg[6] ,
    \value_reg[1]_1 ,
    Q,
    large_error_reg,
    large_error_reg_0,
    get_terminator,
    jumbo_enable,
    large_error_i_4,
    \value_reg[9]_0 ,
    tagged_frame,
    vlan_enable,
    clk_i,
    reset_dcm,
    \value_reg[10]_0 ,
    \value_reg[7] ,
    \value_reg[6]_0 ,
    \value_reg[5] ,
    \value_reg[0] );
  output [6:0]\value_reg[10] ;
  output \value_reg[9] ;
  output \value_reg[11] ;
  output \value_reg[2] ;
  output jumbo_frame0;
  output \value_reg[8] ;
  output \value_reg[4] ;
  output \value_reg[1] ;
  output \value_reg[1]_0 ;
  output length_256_5110;
  output length_512_10230;
  output length_65_1270;
  output padded_frame0;
  output small_error0;
  output length_128_2550;
  output \value_reg[6] ;
  input [0:0]\value_reg[1]_1 ;
  input [2:0]Q;
  input large_error_reg;
  input large_error_reg_0;
  input get_terminator;
  input jumbo_enable;
  input [0:0]large_error_i_4;
  input \value_reg[9]_0 ;
  input tagged_frame;
  input vlan_enable;
  input clk_i;
  input reset_dcm;
  input \value_reg[10]_0 ;
  input \value_reg[7] ;
  input \value_reg[6]_0 ;
  input \value_reg[5] ;
  input \value_reg[0] ;

  wire [2:0]Q;
  wire clk_i;
  wire get_terminator;
  wire jumbo_enable;
  wire jumbo_frame0;
  wire [0:0]large_error_i_4;
  wire large_error_reg;
  wire large_error_reg_0;
  wire length_128_2550;
  wire length_256_5110;
  wire length_512_10230;
  wire length_65_1270;
  wire padded_frame0;
  wire reset_dcm;
  wire small_error0;
  wire tagged_frame;
  wire \value_reg[0] ;
  wire [6:0]\value_reg[10] ;
  wire \value_reg[10]_0 ;
  wire \value_reg[11] ;
  wire \value_reg[1] ;
  wire \value_reg[1]_0 ;
  wire [0:0]\value_reg[1]_1 ;
  wire \value_reg[2] ;
  wire \value_reg[4] ;
  wire \value_reg[5] ;
  wire \value_reg[6] ;
  wire \value_reg[6]_0 ;
  wire \value_reg[7] ;
  wire \value_reg[8] ;
  wire \value_reg[9] ;
  wire \value_reg[9]_0 ;
  wire vlan_enable;

  switch_elements_counter data_counter
       (.Q(Q),
        .clk_i(clk_i),
        .get_terminator(get_terminator),
        .jumbo_enable(jumbo_enable),
        .jumbo_frame0(jumbo_frame0),
        .large_error_i_4_0(large_error_i_4),
        .large_error_reg(large_error_reg),
        .large_error_reg_0(large_error_reg_0),
        .length_128_2550(length_128_2550),
        .length_256_5110(length_256_5110),
        .length_512_10230(length_512_10230),
        .length_65_1270(length_65_1270),
        .padded_frame0(padded_frame0),
        .reset_dcm(reset_dcm),
        .small_error0(small_error0),
        .tagged_frame(tagged_frame),
        .\value_reg[0]_0 (\value_reg[10] [0]),
        .\value_reg[0]_1 (\value_reg[0] ),
        .\value_reg[10]_0 (\value_reg[10] [6]),
        .\value_reg[10]_1 (\value_reg[10]_0 ),
        .\value_reg[11]_0 (\value_reg[11] ),
        .\value_reg[1]_0 (\value_reg[10] [1]),
        .\value_reg[1]_1 (\value_reg[1] ),
        .\value_reg[1]_2 (\value_reg[1]_0 ),
        .\value_reg[1]_3 (\value_reg[1]_1 ),
        .\value_reg[2]_0 (\value_reg[2] ),
        .\value_reg[4]_0 (\value_reg[10] [2]),
        .\value_reg[4]_1 (\value_reg[4] ),
        .\value_reg[5]_0 (\value_reg[10] [3]),
        .\value_reg[5]_1 (\value_reg[5] ),
        .\value_reg[6]_0 (\value_reg[10] [4]),
        .\value_reg[6]_1 (\value_reg[6] ),
        .\value_reg[6]_2 (\value_reg[6]_0 ),
        .\value_reg[7]_0 (\value_reg[10] [5]),
        .\value_reg[7]_1 (\value_reg[7] ),
        .\value_reg[8]_0 (\value_reg[8] ),
        .\value_reg[9]_0 (\value_reg[9] ),
        .\value_reg[9]_1 (\value_reg[9]_0 ),
        .vlan_enable(vlan_enable));
endmodule

(* ORIG_REF_NAME = "rxRSIO" *) 
module switch_elements_rxRSIO
   (AR,
    local_fault,
    remote_fault,
    \FSM_sequential_linkstate_reg[1] ,
    this_cycle,
    D,
    E,
    qvDataOut,
    \qvDataOut_reg[69] ,
    \qvDataOut_reg[62] ,
    get_sfd0,
    \qvDataOut_reg[45] ,
    clk_i,
    Q,
    \rxd32_in_tmp_reg[31]_0 ,
    \rxc4_in_tmp_reg[3]_0 ,
    rst_i,
    recv_rst);
  output [0:0]AR;
  output local_fault;
  output remote_fault;
  output \FSM_sequential_linkstate_reg[1] ;
  output this_cycle;
  output [5:0]D;
  output [0:0]E;
  output [71:0]qvDataOut;
  output [2:0]\qvDataOut_reg[69] ;
  output [7:0]\qvDataOut_reg[62] ;
  output get_sfd0;
  output \qvDataOut_reg[45] ;
  input clk_i;
  input [0:0]Q;
  input [31:0]\rxd32_in_tmp_reg[31]_0 ;
  input [3:0]\rxc4_in_tmp_reg[3]_0 ;
  input rst_i;
  input recv_rst;

  wire [0:0]AR;
  wire [5:0]D;
  wire [0:0]E;
  wire \FSM_sequential_linkstate_reg[1] ;
  wire [71:0]MemDataIn;
  wire [0:0]Q;
  wire clk_i;
  wire get_align_reg;
  wire get_align_reg_i_1_n_0;
  wire get_align_reg_i_2_n_0;
  wire get_align_reg_i_3_n_0;
  wire get_align_reg_i_4_n_0;
  wire get_align_reg_i_5_n_0;
  wire get_align_reg_i_6_n_0;
  wire get_align_reg_i_7_n_0;
  wire get_align_reg_i_8_n_0;
  wire get_align_reg_i_9_n_0;
  wire get_sfd0;
  wire local_fault;
  wire local_fault0;
  wire local_fault3;
  wire local_fault44_in;
  wire local_fault_i_2_n_0;
  wire local_fault_i_3_n_0;
  wire local_fault_i_5_n_0;
  wire local_fault_i_7_n_0;
  wire local_fault_i_8_n_0;
  wire local_fault_i_9_n_0;
  wire p_0_in;
  wire [71:0]qvDataOut;
  wire \qvDataOut_reg[45] ;
  wire [7:0]\qvDataOut_reg[62] ;
  wire [2:0]\qvDataOut_reg[69] ;
  wire \qvWriteCntrl[0]_i_1_n_0 ;
  wire \qvWriteCntrl[1]_i_1_n_0 ;
  wire \qvWriteCntrl_reg_n_0_[0] ;
  wire recv_rst;
  wire remote_fault;
  wire remote_fault0;
  wire rst_i;
  wire [3:0]rxc4_in_tmp_d1;
  wire [3:0]\rxc4_in_tmp_reg[3]_0 ;
  wire \rxc4_in_tmp_reg_n_0_[0] ;
  wire \rxc4_in_tmp_reg_n_0_[1] ;
  wire \rxc4_in_tmp_reg_n_0_[2] ;
  wire \rxc4_in_tmp_reg_n_0_[3] ;
  wire [31:0]rxd32_in_tmp;
  wire [31:0]rxd32_in_tmp_d1;
  wire [31:0]\rxd32_in_tmp_reg[31]_0 ;
  wire \rxd64_in_tmp[31]_i_1_n_0 ;
  wire this_cycle;

  LUT3 #(
    .INIT(8'hFE)) 
    \FSM_sequential_linkstate[0]_i_4 
       (.I0(Q),
        .I1(local_fault),
        .I2(remote_fault),
        .O(\FSM_sequential_linkstate_reg[1] ));
  switch_elements_SwitchAsyncFIFO RealignInst
       (.D(D),
        .E(E),
        .MemDataIn(MemDataIn),
        .Q(\qvWriteCntrl_reg_n_0_[0] ),
        .clk_i(clk_i),
        .get_sfd0(get_sfd0),
        .\qvDataOut_reg[45] (\qvDataOut_reg[45] ),
        .\qvDataOut_reg[62] (\qvDataOut_reg[62] ),
        .\qvDataOut_reg[69] (\qvDataOut_reg[69] ),
        .\qvDataOut_reg[71] (qvDataOut),
        .recv_rst(recv_rst),
        .rst_i(rst_i),
        .rst_i_0(AR),
        .this_cycle(this_cycle));
  LUT6 #(
    .INIT(64'h8000FFFF80008000)) 
    get_align_reg_i_1
       (.I0(\rxc4_in_tmp_reg_n_0_[0] ),
        .I1(rxd32_in_tmp[0]),
        .I2(rxd32_in_tmp[1]),
        .I3(get_align_reg_i_2_n_0),
        .I4(get_align_reg_i_3_n_0),
        .I5(get_align_reg),
        .O(get_align_reg_i_1_n_0));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    get_align_reg_i_2
       (.I0(rxd32_in_tmp[4]),
        .I1(rxd32_in_tmp[5]),
        .I2(rxd32_in_tmp[3]),
        .I3(rxd32_in_tmp[2]),
        .I4(rxd32_in_tmp[7]),
        .I5(rxd32_in_tmp[6]),
        .O(get_align_reg_i_2_n_0));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    get_align_reg_i_3
       (.I0(get_align_reg_i_4_n_0),
        .I1(get_align_reg_i_5_n_0),
        .I2(get_align_reg_i_6_n_0),
        .I3(get_align_reg_i_7_n_0),
        .I4(get_align_reg_i_8_n_0),
        .I5(get_align_reg_i_9_n_0),
        .O(get_align_reg_i_3_n_0));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    get_align_reg_i_4
       (.I0(rxd32_in_tmp[22]),
        .I1(rxd32_in_tmp[23]),
        .I2(rxd32_in_tmp[20]),
        .I3(rxd32_in_tmp[21]),
        .I4(rxd32_in_tmp[25]),
        .I5(rxd32_in_tmp[24]),
        .O(get_align_reg_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    get_align_reg_i_5
       (.I0(rxd32_in_tmp[16]),
        .I1(rxd32_in_tmp[17]),
        .I2(rxd32_in_tmp[14]),
        .I3(rxd32_in_tmp[15]),
        .I4(rxd32_in_tmp[19]),
        .I5(rxd32_in_tmp[18]),
        .O(get_align_reg_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    get_align_reg_i_6
       (.I0(rxd32_in_tmp[1]),
        .I1(rxd32_in_tmp[2]),
        .I2(\rxc4_in_tmp_reg_n_0_[0] ),
        .I3(rxd32_in_tmp[0]),
        .I4(rxd32_in_tmp[4]),
        .I5(rxd32_in_tmp[3]),
        .O(get_align_reg_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    get_align_reg_i_7
       (.I0(rxd32_in_tmp[28]),
        .I1(rxd32_in_tmp[29]),
        .I2(rxd32_in_tmp[26]),
        .I3(rxd32_in_tmp[27]),
        .I4(rxd32_in_tmp[31]),
        .I5(rxd32_in_tmp[30]),
        .O(get_align_reg_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    get_align_reg_i_8
       (.I0(\rxc4_in_tmp_reg_n_0_[3] ),
        .I1(rxd32_in_tmp[5]),
        .I2(\rxc4_in_tmp_reg_n_0_[1] ),
        .I3(\rxc4_in_tmp_reg_n_0_[2] ),
        .I4(rxd32_in_tmp[7]),
        .I5(rxd32_in_tmp[6]),
        .O(get_align_reg_i_8_n_0));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    get_align_reg_i_9
       (.I0(rxd32_in_tmp[10]),
        .I1(rxd32_in_tmp[11]),
        .I2(rxd32_in_tmp[8]),
        .I3(rxd32_in_tmp[9]),
        .I4(rxd32_in_tmp[13]),
        .I5(rxd32_in_tmp[12]),
        .O(get_align_reg_i_9_n_0));
  FDCE #(
    .INIT(1'b0)) 
    get_align_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(get_align_reg_i_1_n_0),
        .Q(get_align_reg));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    local_fault_i_1
       (.I0(\rxd32_in_tmp_reg[31]_0 [30]),
        .I1(\rxd32_in_tmp_reg[31]_0 [31]),
        .I2(local_fault_i_2_n_0),
        .I3(local_fault_i_3_n_0),
        .I4(local_fault44_in),
        .O(local_fault0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    local_fault_i_2
       (.I0(local_fault_i_5_n_0),
        .I1(\rxd32_in_tmp_reg[31]_0 [9]),
        .I2(\rxd32_in_tmp_reg[31]_0 [8]),
        .I3(\rxd32_in_tmp_reg[31]_0 [11]),
        .I4(\rxd32_in_tmp_reg[31]_0 [10]),
        .I5(local_fault3),
        .O(local_fault_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    local_fault_i_3
       (.I0(local_fault_i_7_n_0),
        .I1(\rxd32_in_tmp_reg[31]_0 [23]),
        .I2(\rxd32_in_tmp_reg[31]_0 [22]),
        .I3(\rxd32_in_tmp_reg[31]_0 [21]),
        .I4(\rxd32_in_tmp_reg[31]_0 [20]),
        .I5(local_fault_i_8_n_0),
        .O(local_fault_i_3_n_0));
  LUT5 #(
    .INIT(32'h00200000)) 
    local_fault_i_4
       (.I0(\rxd32_in_tmp_reg[31]_0 [4]),
        .I1(\rxd32_in_tmp_reg[31]_0 [5]),
        .I2(\rxd32_in_tmp_reg[31]_0 [7]),
        .I3(\rxd32_in_tmp_reg[31]_0 [6]),
        .I4(local_fault_i_9_n_0),
        .O(local_fault44_in));
  LUT4 #(
    .INIT(16'h0001)) 
    local_fault_i_5
       (.I0(\rxd32_in_tmp_reg[31]_0 [15]),
        .I1(\rxd32_in_tmp_reg[31]_0 [14]),
        .I2(\rxd32_in_tmp_reg[31]_0 [13]),
        .I3(\rxd32_in_tmp_reg[31]_0 [12]),
        .O(local_fault_i_5_n_0));
  LUT4 #(
    .INIT(16'h0100)) 
    local_fault_i_6
       (.I0(\rxc4_in_tmp_reg[3]_0 [1]),
        .I1(\rxc4_in_tmp_reg[3]_0 [0]),
        .I2(\rxc4_in_tmp_reg[3]_0 [2]),
        .I3(\rxc4_in_tmp_reg[3]_0 [3]),
        .O(local_fault3));
  LUT4 #(
    .INIT(16'h0001)) 
    local_fault_i_7
       (.I0(\rxd32_in_tmp_reg[31]_0 [19]),
        .I1(\rxd32_in_tmp_reg[31]_0 [18]),
        .I2(\rxd32_in_tmp_reg[31]_0 [17]),
        .I3(\rxd32_in_tmp_reg[31]_0 [16]),
        .O(local_fault_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    local_fault_i_8
       (.I0(\rxd32_in_tmp_reg[31]_0 [28]),
        .I1(\rxd32_in_tmp_reg[31]_0 [29]),
        .I2(\rxd32_in_tmp_reg[31]_0 [27]),
        .I3(\rxd32_in_tmp_reg[31]_0 [26]),
        .I4(\rxd32_in_tmp_reg[31]_0 [24]),
        .I5(\rxd32_in_tmp_reg[31]_0 [25]),
        .O(local_fault_i_8_n_0));
  LUT4 #(
    .INIT(16'h0400)) 
    local_fault_i_9
       (.I0(\rxd32_in_tmp_reg[31]_0 [0]),
        .I1(\rxd32_in_tmp_reg[31]_0 [1]),
        .I2(\rxd32_in_tmp_reg[31]_0 [2]),
        .I3(\rxd32_in_tmp_reg[31]_0 [3]),
        .O(local_fault_i_9_n_0));
  FDCE #(
    .INIT(1'b0)) 
    local_fault_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(local_fault0),
        .Q(local_fault));
  LUT2 #(
    .INIT(4'hB)) 
    \qvWriteCntrl[0]_i_1 
       (.I0(p_0_in),
        .I1(get_align_reg),
        .O(\qvWriteCntrl[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \qvWriteCntrl[1]_i_1 
       (.I0(\qvWriteCntrl_reg_n_0_[0] ),
        .I1(get_align_reg),
        .O(\qvWriteCntrl[1]_i_1_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \qvWriteCntrl_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\qvWriteCntrl[0]_i_1_n_0 ),
        .PRE(AR),
        .Q(\qvWriteCntrl_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \qvWriteCntrl_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\qvWriteCntrl[1]_i_1_n_0 ),
        .Q(p_0_in));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    remote_fault_i_1
       (.I0(\rxd32_in_tmp_reg[31]_0 [31]),
        .I1(\rxd32_in_tmp_reg[31]_0 [30]),
        .I2(local_fault_i_2_n_0),
        .I3(local_fault_i_3_n_0),
        .I4(local_fault44_in),
        .O(remote_fault0));
  FDCE #(
    .INIT(1'b0)) 
    remote_fault_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(remote_fault0),
        .Q(remote_fault));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg_n_0_[0] ),
        .Q(rxc4_in_tmp_d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg_n_0_[1] ),
        .Q(rxc4_in_tmp_d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg_n_0_[2] ),
        .Q(rxc4_in_tmp_d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg_n_0_[3] ),
        .Q(rxc4_in_tmp_d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg[3]_0 [0]),
        .Q(\rxc4_in_tmp_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg[3]_0 [1]),
        .Q(\rxc4_in_tmp_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg[3]_0 [2]),
        .Q(\rxc4_in_tmp_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \rxc4_in_tmp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxc4_in_tmp_reg[3]_0 [3]),
        .Q(\rxc4_in_tmp_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[0] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[0]),
        .Q(MemDataIn[64]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[1] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[1]),
        .Q(MemDataIn[65]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[2] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[2]),
        .Q(MemDataIn[66]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[3] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[3]),
        .Q(MemDataIn[67]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[4] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[0]),
        .Q(MemDataIn[68]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[5] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[1]),
        .Q(MemDataIn[69]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[6] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[2]),
        .Q(MemDataIn[70]));
  FDCE #(
    .INIT(1'b0)) 
    \rxc8_in_tmp_reg[7] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxc4_in_tmp_d1[3]),
        .Q(MemDataIn[71]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[0]),
        .Q(rxd32_in_tmp_d1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[10]),
        .Q(rxd32_in_tmp_d1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[11]),
        .Q(rxd32_in_tmp_d1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[12]),
        .Q(rxd32_in_tmp_d1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[13]),
        .Q(rxd32_in_tmp_d1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[14]),
        .Q(rxd32_in_tmp_d1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[15]),
        .Q(rxd32_in_tmp_d1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[16]),
        .Q(rxd32_in_tmp_d1[16]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[17]),
        .Q(rxd32_in_tmp_d1[17]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[18]),
        .Q(rxd32_in_tmp_d1[18]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[19]),
        .Q(rxd32_in_tmp_d1[19]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[1]),
        .Q(rxd32_in_tmp_d1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[20]),
        .Q(rxd32_in_tmp_d1[20]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[21]),
        .Q(rxd32_in_tmp_d1[21]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[22]),
        .Q(rxd32_in_tmp_d1[22]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[23]),
        .Q(rxd32_in_tmp_d1[23]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[24]),
        .Q(rxd32_in_tmp_d1[24]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[25]),
        .Q(rxd32_in_tmp_d1[25]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[26]),
        .Q(rxd32_in_tmp_d1[26]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[27]),
        .Q(rxd32_in_tmp_d1[27]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[28]),
        .Q(rxd32_in_tmp_d1[28]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[29]),
        .Q(rxd32_in_tmp_d1[29]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[2]),
        .Q(rxd32_in_tmp_d1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[30]),
        .Q(rxd32_in_tmp_d1[30]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[31]),
        .Q(rxd32_in_tmp_d1[31]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[3]),
        .Q(rxd32_in_tmp_d1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[4]),
        .Q(rxd32_in_tmp_d1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[5]),
        .Q(rxd32_in_tmp_d1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[6]),
        .Q(rxd32_in_tmp_d1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[7]),
        .Q(rxd32_in_tmp_d1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[8]),
        .Q(rxd32_in_tmp_d1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_d1_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(rxd32_in_tmp[9]),
        .Q(rxd32_in_tmp_d1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [0]),
        .Q(rxd32_in_tmp[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [10]),
        .Q(rxd32_in_tmp[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [11]),
        .Q(rxd32_in_tmp[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [12]),
        .Q(rxd32_in_tmp[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [13]),
        .Q(rxd32_in_tmp[13]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [14]),
        .Q(rxd32_in_tmp[14]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [15]),
        .Q(rxd32_in_tmp[15]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [16]),
        .Q(rxd32_in_tmp[16]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [17]),
        .Q(rxd32_in_tmp[17]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [18]),
        .Q(rxd32_in_tmp[18]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [19]),
        .Q(rxd32_in_tmp[19]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [1]),
        .Q(rxd32_in_tmp[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [20]),
        .Q(rxd32_in_tmp[20]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [21]),
        .Q(rxd32_in_tmp[21]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [22]),
        .Q(rxd32_in_tmp[22]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [23]),
        .Q(rxd32_in_tmp[23]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [24]),
        .Q(rxd32_in_tmp[24]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [25]),
        .Q(rxd32_in_tmp[25]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [26]),
        .Q(rxd32_in_tmp[26]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [27]),
        .Q(rxd32_in_tmp[27]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [28]),
        .Q(rxd32_in_tmp[28]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [29]),
        .Q(rxd32_in_tmp[29]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [2]),
        .Q(rxd32_in_tmp[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [30]),
        .Q(rxd32_in_tmp[30]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [31]),
        .Q(rxd32_in_tmp[31]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [3]),
        .Q(rxd32_in_tmp[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [4]),
        .Q(rxd32_in_tmp[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [5]),
        .Q(rxd32_in_tmp[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [6]),
        .Q(rxd32_in_tmp[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [7]),
        .Q(rxd32_in_tmp[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [8]),
        .Q(rxd32_in_tmp[8]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd32_in_tmp_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(AR),
        .D(\rxd32_in_tmp_reg[31]_0 [9]),
        .Q(rxd32_in_tmp[9]));
  LUT1 #(
    .INIT(2'h1)) 
    \rxd64_in_tmp[31]_i_1 
       (.I0(p_0_in),
        .O(\rxd64_in_tmp[31]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[0] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[0]),
        .Q(MemDataIn[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[10] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[10]),
        .Q(MemDataIn[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[11] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[11]),
        .Q(MemDataIn[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[12] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[12]),
        .Q(MemDataIn[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[13] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[13]),
        .Q(MemDataIn[13]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[14] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[14]),
        .Q(MemDataIn[14]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[15] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[15]),
        .Q(MemDataIn[15]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[16] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[16]),
        .Q(MemDataIn[16]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[17] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[17]),
        .Q(MemDataIn[17]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[18] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[18]),
        .Q(MemDataIn[18]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[19] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[19]),
        .Q(MemDataIn[19]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[1] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[1]),
        .Q(MemDataIn[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[20] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[20]),
        .Q(MemDataIn[20]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[21] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[21]),
        .Q(MemDataIn[21]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[22] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[22]),
        .Q(MemDataIn[22]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[23] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[23]),
        .Q(MemDataIn[23]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[24] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[24]),
        .Q(MemDataIn[24]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[25] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[25]),
        .Q(MemDataIn[25]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[26] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[26]),
        .Q(MemDataIn[26]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[27] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[27]),
        .Q(MemDataIn[27]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[28] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[28]),
        .Q(MemDataIn[28]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[29] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[29]),
        .Q(MemDataIn[29]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[2] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[2]),
        .Q(MemDataIn[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[30] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[30]),
        .Q(MemDataIn[30]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[31] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[31]),
        .Q(MemDataIn[31]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[32] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[0]),
        .Q(MemDataIn[32]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[33] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[1]),
        .Q(MemDataIn[33]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[34] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[2]),
        .Q(MemDataIn[34]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[35] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[3]),
        .Q(MemDataIn[35]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[36] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[4]),
        .Q(MemDataIn[36]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[37] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[5]),
        .Q(MemDataIn[37]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[38] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[6]),
        .Q(MemDataIn[38]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[39] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[7]),
        .Q(MemDataIn[39]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[3] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[3]),
        .Q(MemDataIn[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[40] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[8]),
        .Q(MemDataIn[40]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[41] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[9]),
        .Q(MemDataIn[41]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[42] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[10]),
        .Q(MemDataIn[42]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[43] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[11]),
        .Q(MemDataIn[43]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[44] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[12]),
        .Q(MemDataIn[44]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[45] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[13]),
        .Q(MemDataIn[45]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[46] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[14]),
        .Q(MemDataIn[46]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[47] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[15]),
        .Q(MemDataIn[47]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[48] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[16]),
        .Q(MemDataIn[48]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[49] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[17]),
        .Q(MemDataIn[49]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[4] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[4]),
        .Q(MemDataIn[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[50] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[18]),
        .Q(MemDataIn[50]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[51] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[19]),
        .Q(MemDataIn[51]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[52] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[20]),
        .Q(MemDataIn[52]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[53] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[21]),
        .Q(MemDataIn[53]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[54] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[22]),
        .Q(MemDataIn[54]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[55] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[23]),
        .Q(MemDataIn[55]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[56] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[24]),
        .Q(MemDataIn[56]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[57] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[25]),
        .Q(MemDataIn[57]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[58] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[26]),
        .Q(MemDataIn[58]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[59] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[27]),
        .Q(MemDataIn[59]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[5] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[5]),
        .Q(MemDataIn[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[60] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[28]),
        .Q(MemDataIn[60]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[61] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[29]),
        .Q(MemDataIn[61]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[62] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[30]),
        .Q(MemDataIn[62]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[63] 
       (.C(clk_i),
        .CE(p_0_in),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[31]),
        .Q(MemDataIn[63]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[6] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[6]),
        .Q(MemDataIn[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[7] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[7]),
        .Q(MemDataIn[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[8] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[8]),
        .Q(MemDataIn[8]));
  FDCE #(
    .INIT(1'b0)) 
    \rxd64_in_tmp_reg[9] 
       (.C(clk_i),
        .CE(\rxd64_in_tmp[31]_i_1_n_0 ),
        .CLR(AR),
        .D(rxd32_in_tmp_d1[9]),
        .Q(MemDataIn[9]));
endmodule

(* ORIG_REF_NAME = "rxRSLayer" *) 
module switch_elements_rxRSLayer
   (reset_dcm,
    this_cycle,
    D,
    E,
    Q,
    \link_fault_reg[1] ,
    \qvDataOut_reg[69] ,
    \qvDataOut_reg[62] ,
    get_sfd0,
    \qvDataOut_reg[45] ,
    clk_i,
    rxclk_180,
    \rxd32_in_tmp_reg[31] ,
    \rxc4_in_tmp_reg[3] ,
    rst_i,
    recv_rst);
  output reset_dcm;
  output this_cycle;
  output [5:0]D;
  output [0:0]E;
  output [71:0]Q;
  output [1:0]\link_fault_reg[1] ;
  output [2:0]\qvDataOut_reg[69] ;
  output [7:0]\qvDataOut_reg[62] ;
  output get_sfd0;
  output \qvDataOut_reg[45] ;
  input clk_i;
  input rxclk_180;
  input [31:0]\rxd32_in_tmp_reg[31] ;
  input [3:0]\rxc4_in_tmp_reg[3] ;
  input rst_i;
  input recv_rst;

  wire [5:0]D;
  wire [0:0]E;
  wire [71:0]Q;
  wire clk_i;
  wire datapath_n_3;
  wire get_sfd0;
  wire [1:0]\link_fault_reg[1] ;
  wire [1:1]linkstate;
  wire local_fault;
  wire \qvDataOut_reg[45] ;
  wire [7:0]\qvDataOut_reg[62] ;
  wire [2:0]\qvDataOut_reg[69] ;
  wire recv_rst;
  wire remote_fault;
  wire reset_dcm;
  wire rst_i;
  wire [3:0]\rxc4_in_tmp_reg[3] ;
  wire rxclk_180;
  wire [31:0]\rxd32_in_tmp_reg[31] ;
  wire this_cycle;

  switch_elements_rxRSIO datapath
       (.AR(reset_dcm),
        .D(D),
        .E(E),
        .\FSM_sequential_linkstate_reg[1] (datapath_n_3),
        .Q(linkstate),
        .clk_i(clk_i),
        .get_sfd0(get_sfd0),
        .local_fault(local_fault),
        .qvDataOut(Q),
        .\qvDataOut_reg[45] (\qvDataOut_reg[45] ),
        .\qvDataOut_reg[62] (\qvDataOut_reg[62] ),
        .\qvDataOut_reg[69] (\qvDataOut_reg[69] ),
        .recv_rst(recv_rst),
        .remote_fault(remote_fault),
        .rst_i(rst_i),
        .\rxc4_in_tmp_reg[3]_0 (\rxc4_in_tmp_reg[3] ),
        .\rxd32_in_tmp_reg[31]_0 (\rxd32_in_tmp_reg[31] ),
        .this_cycle(this_cycle));
  switch_elements_rxLinkFaultState statemachine
       (.AR(reset_dcm),
        .\FSM_sequential_linkstate_reg[0]_0 (datapath_n_3),
        .Q(linkstate),
        .\link_fault_reg[1]_0 (\link_fault_reg[1] ),
        .local_fault(local_fault),
        .remote_fault(remote_fault),
        .rxclk_180(rxclk_180));
endmodule

(* ORIG_REF_NAME = "rxReceiveEngine" *) 
module switch_elements_rxReceiveEngine
   (in0,
    rx_bad_frame,
    rx_good_frame,
    rxCfgofRS,
    Q,
    rx_data_valid,
    rx_data,
    clk_i,
    rxclk_180,
    rst_i,
    D,
    \rxc4_in_tmp_reg[3] ,
    \cfgRxRegData_reg[52]_0 );
  output [13:0]in0;
  output rx_bad_frame;
  output rx_good_frame;
  output [2:0]rxCfgofRS;
  output [1:0]Q;
  output [7:0]rx_data_valid;
  output [63:0]rx_data;
  input clk_i;
  input rxclk_180;
  input rst_i;
  input [31:0]D;
  input [3:0]\rxc4_in_tmp_reg[3] ;
  input [4:0]\cfgRxRegData_reg[52]_0 ;

  wire [31:0]D;
  wire [1:0]Q;
  wire bad_frame_get;
  wire bad_frame_get0;
  wire broad_valid;
  wire [1:0]bytes_cnt;
  wire [4:0]\cfgRxRegData_reg[52]_0 ;
  wire \cfgRxRegData_reg_n_0_[48] ;
  wire \cfgRxRegData_reg_n_0_[49] ;
  wire \cfgRxRegData_reg_n_0_[50] ;
  wire \cfgRxRegData_reg_n_0_[51] ;
  wire \cfgRxRegData_reg_n_0_[52] ;
  wire check_reset;
  wire clk_i;
  wire counters_n_11;
  wire counters_n_12;
  wire counters_n_13;
  wire counters_n_14;
  wire counters_n_21;
  wire counters_n_7;
  wire counters_n_8;
  wire counters_n_9;
  wire \crc64/nextCRC32_D64_return0 ;
  wire \crc64/nextCRC32_D64_return0100_out ;
  wire \crc64/nextCRC32_D64_return0102_out ;
  wire \crc64/nextCRC32_D64_return0104_out ;
  wire \crc64/nextCRC32_D64_return0106_out ;
  wire \crc64/nextCRC32_D64_return0108_out ;
  wire \crc64/nextCRC32_D64_return0109_out ;
  wire \crc64/nextCRC32_D64_return0110_out ;
  wire \crc64/nextCRC32_D64_return0112_out ;
  wire \crc64/nextCRC32_D64_return0114_out ;
  wire \crc64/nextCRC32_D64_return0116_out ;
  wire \crc64/nextCRC32_D64_return0118_out ;
  wire \crc64/nextCRC32_D64_return0120_out ;
  wire \crc64/nextCRC32_D64_return0122_out ;
  wire \crc64/nextCRC32_D64_return0124_out ;
  wire \crc64/nextCRC32_D64_return0126_out ;
  wire \crc64/nextCRC32_D64_return0128_out ;
  wire \crc64/nextCRC32_D64_return0130_out ;
  wire \crc64/nextCRC32_D64_return0132_out ;
  wire \crc64/nextCRC32_D64_return0136_out ;
  wire \crc64/nextCRC32_D64_return0138_out ;
  wire \crc64/nextCRC32_D64_return056_out ;
  wire \crc64/nextCRC32_D64_return068_out ;
  wire \crc64/nextCRC32_D64_return075_out ;
  wire \crc64/nextCRC32_D64_return080_out ;
  wire \crc64/nextCRC32_D64_return086_out ;
  wire \crc64/nextCRC32_D64_return091_out ;
  wire \crc64/nextCRC32_D64_return093_out ;
  wire \crc64/nextCRC32_D64_return094_out ;
  wire \crc64/nextCRC32_D64_return096_out ;
  wire \crc64/nextCRC32_D64_return098_out ;
  wire crc_64_en;
  wire crc_check_invalid;
  wire [31:0]crc_from_64;
  wire crcmodule_n_4;
  wire crcmodule_n_40;
  wire crcmodule_n_41;
  wire crcmodule_n_42;
  wire crcmodule_n_43;
  wire crcmodule_n_44;
  wire crcmodule_n_45;
  wire crcmodule_n_46;
  wire crcmodule_n_47;
  wire crcmodule_n_48;
  wire crcmodule_n_49;
  wire crcmodule_n_5;
  wire crcmodule_n_50;
  wire crcmodule_n_51;
  wire crcmodule_n_52;
  wire crcmodule_n_53;
  wire crcmodule_n_54;
  wire crcmodule_n_55;
  wire crcmodule_n_56;
  wire crcmodule_n_57;
  wire crcmodule_n_58;
  wire crcmodule_n_59;
  wire crcmodule_n_60;
  wire crcmodule_n_61;
  wire crcmodule_n_62;
  wire crcmodule_n_63;
  wire crcmodule_n_64;
  wire crcmodule_n_65;
  wire crcmodule_n_66;
  wire crcmodule_n_67;
  wire crcmodule_n_68;
  wire crcmodule_n_69;
  wire crcmodule_n_70;
  wire crcmodule_n_71;
  wire crcmodule_n_72;
  wire crcmodule_n_73;
  wire crcmodule_n_74;
  wire crcmodule_n_75;
  wire crcmodule_n_76;
  wire crcmodule_n_77;
  wire crcmodule_n_78;
  wire crcmodule_n_79;
  wire crcmodule_n_9;
  wire datapath_main_n_112;
  wire datapath_main_n_113;
  wire datapath_main_n_114;
  wire datapath_main_n_115;
  wire datapath_main_n_116;
  wire datapath_main_n_117;
  wire datapath_main_n_118;
  wire datapath_main_n_119;
  wire datapath_main_n_120;
  wire datapath_main_n_121;
  wire datapath_main_n_194;
  wire datapath_main_n_195;
  wire datapath_main_n_73;
  wire datapath_main_n_74;
  wire datapath_main_n_75;
  wire datapath_main_n_79;
  wire datapath_main_n_80;
  wire do_crc_check;
  wire [0:0]fifo_state;
  wire [10:0]frame_cnt;
  wire get_error_code;
  wire get_sfd;
  wire get_sfd0;
  wire get_terminator;
  wire get_terminator_d1;
  wire get_terminator_d2;
  wire get_terminator_d3;
  wire good_frame_get;
  wire [13:0]in0;
  wire inband_fcs;
  wire jumbo_enable;
  wire jumbo_frame;
  wire jumbo_frame0;
  wire large_error;
  wire lenchecker_n_11;
  wire lenchecker_n_13;
  wire lenchecker_n_8;
  wire lenchecker_n_9;
  wire length_128_255;
  wire length_128_2550;
  wire length_256_511;
  wire length_256_5110;
  wire length_512_1023;
  wire length_512_10230;
  wire length_65_127;
  wire length_65_1270;
  wire [2:2]location_reg;
  wire multi_valid;
  wire [1:1]p_0_in;
  wire [7:0]p_16_out;
  wire padded_frame;
  wire padded_frame0;
  wire receiving;
  wire recv_enable;
  wire recv_rst;
  wire reset_dcm;
  wire rst_i;
  wire [2:0]rxCfgofRS;
  wire rxStatRegPlus_tmp0;
  wire rxStatRegPlus_tmp00_out;
  wire rxStatRegPlus_tmp01_out;
  wire rxStatRegPlus_tmp02_out;
  wire rxStatRegPlus_tmp03_out;
  wire rxStatRegPlus_tmp04_out;
  wire rxStatRegPlus_tmp05_out;
  wire rxStatRegPlus_tmp08_out;
  wire rxStatRegPlus_tmp09_out;
  wire rx_bad_frame;
  wire [63:0]rx_data;
  wire [7:0]rx_data_valid;
  wire rx_good_frame;
  wire rx_rs_n_2;
  wire rx_rs_n_3;
  wire rx_rs_n_4;
  wire rx_rs_n_5;
  wire rx_rs_n_6;
  wire rx_rs_n_7;
  wire rx_rs_n_83;
  wire rx_rs_n_84;
  wire rx_rs_n_85;
  wire rx_rs_n_95;
  wire [3:0]\rxc4_in_tmp_reg[3] ;
  wire [7:0]rxc8;
  wire rxclk_180;
  wire [63:0]rxd64;
  wire [63:0]rxd64_d3;
  wire small_error;
  wire small_error0;
  wire start_da;
  wire start_lt;
  wire statemachine_n_13;
  wire statemachine_n_14;
  wire statemachine_n_19;
  wire statemachine_n_20;
  wire statemachine_n_21;
  wire statemachine_n_22;
  wire statemachine_n_23;
  wire statemachine_n_24;
  wire statemachine_n_25;
  wire tagged_frame;
  wire [2:0]terminator_location;
  wire terminator_location0;
  wire this_cycle;
  wire vlan_enable;
  wire wait_crc_check;

  FDCE #(
    .INIT(1'b0)) 
    \cfgRxRegData_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg[52]_0 [0]),
        .Q(\cfgRxRegData_reg_n_0_[48] ));
  FDCE #(
    .INIT(1'b0)) 
    \cfgRxRegData_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg[52]_0 [1]),
        .Q(\cfgRxRegData_reg_n_0_[49] ));
  FDCE #(
    .INIT(1'b0)) 
    \cfgRxRegData_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg[52]_0 [2]),
        .Q(\cfgRxRegData_reg_n_0_[50] ));
  FDCE #(
    .INIT(1'b0)) 
    \cfgRxRegData_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg[52]_0 [3]),
        .Q(\cfgRxRegData_reg_n_0_[51] ));
  FDCE #(
    .INIT(1'b0)) 
    \cfgRxRegData_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg[52]_0 [4]),
        .Q(\cfgRxRegData_reg_n_0_[52] ));
  switch_elements_rxNumCounter counters
       (.Q({statemachine_n_14,start_lt,start_da}),
        .clk_i(clk_i),
        .get_terminator(get_terminator),
        .jumbo_enable(jumbo_enable),
        .jumbo_frame0(jumbo_frame0),
        .large_error_i_4(location_reg),
        .large_error_reg(lenchecker_n_13),
        .large_error_reg_0(lenchecker_n_11),
        .length_128_2550(length_128_2550),
        .length_256_5110(length_256_5110),
        .length_512_10230(length_512_10230),
        .length_65_1270(length_65_1270),
        .padded_frame0(padded_frame0),
        .reset_dcm(reset_dcm),
        .small_error0(small_error0),
        .tagged_frame(tagged_frame),
        .\value_reg[0] (statemachine_n_21),
        .\value_reg[10] ({frame_cnt[10],frame_cnt[7:4],frame_cnt[1:0]}),
        .\value_reg[10]_0 (statemachine_n_25),
        .\value_reg[11] (counters_n_8),
        .\value_reg[1] (counters_n_13),
        .\value_reg[1]_0 (counters_n_14),
        .\value_reg[1]_1 (p_0_in),
        .\value_reg[2] (counters_n_9),
        .\value_reg[4] (counters_n_12),
        .\value_reg[5] (statemachine_n_22),
        .\value_reg[6] (counters_n_21),
        .\value_reg[6]_0 (statemachine_n_23),
        .\value_reg[7] (statemachine_n_24),
        .\value_reg[8] (counters_n_11),
        .\value_reg[9] (counters_n_7),
        .\value_reg[9]_0 (statemachine_n_19),
        .vlan_enable(vlan_enable));
  switch_elements_rxCRC crcmodule
       (.\CRC_OUT_reg[0] (crcmodule_n_74),
        .\CRC_OUT_reg[10] (crcmodule_n_64),
        .\CRC_OUT_reg[11] (crcmodule_n_44),
        .\CRC_OUT_reg[14] (crcmodule_n_47),
        .\CRC_OUT_reg[15] (crcmodule_n_52),
        .\CRC_OUT_reg[15]_0 (crcmodule_n_56),
        .\CRC_OUT_reg[15]_1 (crcmodule_n_59),
        .\CRC_OUT_reg[16] (crcmodule_n_76),
        .\CRC_OUT_reg[17] (crcmodule_n_49),
        .\CRC_OUT_reg[18] (crcmodule_n_45),
        .\CRC_OUT_reg[19] (crcmodule_n_65),
        .\CRC_OUT_reg[1] (datapath_main_n_112),
        .\CRC_OUT_reg[20] (crcmodule_n_71),
        .\CRC_OUT_reg[22] (crcmodule_n_70),
        .\CRC_OUT_reg[22]_0 (datapath_main_n_117),
        .\CRC_OUT_reg[22]_1 (datapath_main_n_115),
        .\CRC_OUT_reg[23] (crcmodule_n_79),
        .\CRC_OUT_reg[24] (datapath_main_n_116),
        .\CRC_OUT_reg[24]_0 (datapath_main_n_113),
        .\CRC_OUT_reg[24]_1 (datapath_main_n_118),
        .\CRC_OUT_reg[25] (crcmodule_n_42),
        .\CRC_OUT_reg[26] (crcmodule_n_53),
        .\CRC_OUT_reg[26]_0 (crcmodule_n_61),
        .\CRC_OUT_reg[27] (crcmodule_n_50),
        .\CRC_OUT_reg[28] (crcmodule_n_55),
        .\CRC_OUT_reg[28]_0 (crcmodule_n_57),
        .\CRC_OUT_reg[28]_1 (crcmodule_n_58),
        .\CRC_OUT_reg[29] (crcmodule_n_40),
        .\CRC_OUT_reg[29]_0 (crcmodule_n_41),
        .\CRC_OUT_reg[29]_1 (crcmodule_n_72),
        .\CRC_OUT_reg[29]_2 (datapath_main_n_119),
        .\CRC_OUT_reg[29]_3 (datapath_main_n_120),
        .\CRC_OUT_reg[29]_4 (datapath_main_n_114),
        .\CRC_OUT_reg[2] (crcmodule_n_60),
        .\CRC_OUT_reg[30] (crcmodule_n_54),
        .\CRC_OUT_reg[30]_0 (crcmodule_n_66),
        .\CRC_OUT_reg[30]_1 (crcmodule_n_67),
        .\CRC_OUT_reg[31] ({crc_from_64[31:30],crc_from_64[28:10],crc_from_64[8:0]}),
        .\CRC_OUT_reg[31]_0 (crcmodule_n_75),
        .\CRC_OUT_reg[31]_1 ({\crc64/nextCRC32_D64_return0138_out ,\crc64/nextCRC32_D64_return0136_out ,\crc64/nextCRC32_D64_return0132_out ,\crc64/nextCRC32_D64_return0130_out ,\crc64/nextCRC32_D64_return0128_out ,\crc64/nextCRC32_D64_return0126_out ,\crc64/nextCRC32_D64_return0124_out ,\crc64/nextCRC32_D64_return0122_out ,\crc64/nextCRC32_D64_return0120_out ,\crc64/nextCRC32_D64_return0118_out ,\crc64/nextCRC32_D64_return0116_out ,\crc64/nextCRC32_D64_return0114_out ,\crc64/nextCRC32_D64_return0112_out ,\crc64/nextCRC32_D64_return0110_out ,\crc64/nextCRC32_D64_return0109_out ,\crc64/nextCRC32_D64_return0108_out ,\crc64/nextCRC32_D64_return0106_out ,\crc64/nextCRC32_D64_return0104_out ,\crc64/nextCRC32_D64_return0102_out ,\crc64/nextCRC32_D64_return0100_out ,\crc64/nextCRC32_D64_return098_out ,\crc64/nextCRC32_D64_return096_out ,\crc64/nextCRC32_D64_return094_out ,\crc64/nextCRC32_D64_return093_out ,\crc64/nextCRC32_D64_return091_out ,\crc64/nextCRC32_D64_return086_out ,\crc64/nextCRC32_D64_return080_out ,\crc64/nextCRC32_D64_return075_out ,\crc64/nextCRC32_D64_return068_out ,\crc64/nextCRC32_D64_return056_out ,\crc64/nextCRC32_D64_return0 }),
        .\CRC_OUT_reg[3] (crcmodule_n_69),
        .\CRC_OUT_reg[3]_0 (crcmodule_n_73),
        .\CRC_OUT_reg[6] (datapath_main_n_121),
        .\CRC_OUT_reg[7] (crcmodule_n_48),
        .\CRC_OUT_reg[9] (crcmodule_n_68),
        .\CRC_OUT_reg[9]_0 (crcmodule_n_78),
        .D(crc_check_invalid),
        .E(datapath_main_n_73),
        .Q(statemachine_n_13),
        .SS(datapath_main_n_80),
        .\bytes_cnt_reg[1]_0 (bytes_cnt),
        .\bytes_cnt_reg[1]_1 ({datapath_main_n_74,datapath_main_n_75}),
        .\bytes_cnt_reg[2]_0 (crcmodule_n_9),
        .\bytes_cnt_reg[2]_1 (terminator_location[2]),
        .clk_i(clk_i),
        .crc_64_en(crc_64_en),
        .crc_8_en_reg_0(crcmodule_n_4),
        .do_crc_check(do_crc_check),
        .do_crc_check_reg_0(datapath_main_n_79),
        .get_terminator(get_terminator),
        .get_terminator_d1(get_terminator_d1),
        .get_terminator_d2(get_terminator_d2),
        .get_terminator_d3(get_terminator_d3),
        .large_error(large_error),
        .reset_dcm(reset_dcm),
        .rxd64_d3(rxd64_d3),
        .\rxd64_d3_reg[2] (crcmodule_n_62),
        .\rxd64_d3_reg[33] (crcmodule_n_63),
        .\rxd64_d3_reg[37] (crcmodule_n_43),
        .\rxd64_d3_reg[37]_0 (crcmodule_n_77),
        .\rxd64_d3_reg[48] (crcmodule_n_46),
        .\rxd64_d3_reg[54] (crcmodule_n_51),
        .small_error(small_error),
        .small_error_reg(crcmodule_n_5),
        .wait_crc_check(wait_crc_check));
  switch_elements_rxDAchecker dachecker
       (.broad_valid(broad_valid),
        .broad_valid_reg_0(datapath_main_n_194),
        .clk_i(clk_i),
        .multi_valid(multi_valid),
        .multi_valid_reg_0(datapath_main_n_195),
        .reset_dcm(reset_dcm));
  switch_elements_rxDataPath datapath_main
       (.\CRC_OUT_reg[10] (crcmodule_n_67),
        .\CRC_OUT_reg[11] (crcmodule_n_61),
        .\CRC_OUT_reg[11]_0 (crcmodule_n_45),
        .\CRC_OUT_reg[12] (crcmodule_n_63),
        .\CRC_OUT_reg[13] (crcmodule_n_70),
        .\CRC_OUT_reg[13]_0 (crcmodule_n_42),
        .\CRC_OUT_reg[14] (crcmodule_n_77),
        .\CRC_OUT_reg[14]_0 (crcmodule_n_75),
        .\CRC_OUT_reg[15] (crcmodule_n_79),
        .\CRC_OUT_reg[15]_0 (crcmodule_n_71),
        .\CRC_OUT_reg[16] (crcmodule_n_56),
        .\CRC_OUT_reg[17] (crcmodule_n_49),
        .\CRC_OUT_reg[18] (datapath_main_n_118),
        .\CRC_OUT_reg[18]_0 (crcmodule_n_46),
        .\CRC_OUT_reg[18]_1 (crcmodule_n_76),
        .\CRC_OUT_reg[18]_2 (crcmodule_n_60),
        .\CRC_OUT_reg[1] ({crc_from_64[31:30],crc_from_64[28:10],crc_from_64[8:0]}),
        .\CRC_OUT_reg[1]_0 (crcmodule_n_51),
        .\CRC_OUT_reg[20] (crcmodule_n_48),
        .\CRC_OUT_reg[22] (crcmodule_n_57),
        .\CRC_OUT_reg[22]_0 (crcmodule_n_53),
        .\CRC_OUT_reg[23] (crcmodule_n_52),
        .\CRC_OUT_reg[24] (crcmodule_n_40),
        .\CRC_OUT_reg[24]_0 (crcmodule_n_73),
        .\CRC_OUT_reg[25] (crcmodule_n_41),
        .\CRC_OUT_reg[26] (crcmodule_n_59),
        .\CRC_OUT_reg[27] ({\crc64/nextCRC32_D64_return0138_out ,\crc64/nextCRC32_D64_return0136_out ,\crc64/nextCRC32_D64_return0132_out ,\crc64/nextCRC32_D64_return0130_out ,\crc64/nextCRC32_D64_return0128_out ,\crc64/nextCRC32_D64_return0126_out ,\crc64/nextCRC32_D64_return0124_out ,\crc64/nextCRC32_D64_return0122_out ,\crc64/nextCRC32_D64_return0120_out ,\crc64/nextCRC32_D64_return0118_out ,\crc64/nextCRC32_D64_return0116_out ,\crc64/nextCRC32_D64_return0114_out ,\crc64/nextCRC32_D64_return0112_out ,\crc64/nextCRC32_D64_return0110_out ,\crc64/nextCRC32_D64_return0109_out ,\crc64/nextCRC32_D64_return0108_out ,\crc64/nextCRC32_D64_return0106_out ,\crc64/nextCRC32_D64_return0104_out ,\crc64/nextCRC32_D64_return0102_out ,\crc64/nextCRC32_D64_return0100_out ,\crc64/nextCRC32_D64_return098_out ,\crc64/nextCRC32_D64_return096_out ,\crc64/nextCRC32_D64_return094_out ,\crc64/nextCRC32_D64_return093_out ,\crc64/nextCRC32_D64_return091_out ,\crc64/nextCRC32_D64_return086_out ,\crc64/nextCRC32_D64_return080_out ,\crc64/nextCRC32_D64_return075_out ,\crc64/nextCRC32_D64_return068_out ,\crc64/nextCRC32_D64_return056_out ,\crc64/nextCRC32_D64_return0 }),
        .\CRC_OUT_reg[28] (crcmodule_n_43),
        .\CRC_OUT_reg[28]_0 (crcmodule_n_66),
        .\CRC_OUT_reg[30] (crcmodule_n_69),
        .\CRC_OUT_reg[31] (crcmodule_n_58),
        .\CRC_OUT_reg[4] (crcmodule_n_50),
        .\CRC_OUT_reg[5] (datapath_main_n_116),
        .\CRC_OUT_reg[5]_0 (crcmodule_n_78),
        .\CRC_OUT_reg[5]_1 (crcmodule_n_62),
        .\CRC_OUT_reg[6] (datapath_main_n_115),
        .\CRC_OUT_reg[6]_0 (crcmodule_n_54),
        .\CRC_OUT_reg[6]_1 (crcmodule_n_44),
        .\CRC_OUT_reg[8] (crcmodule_n_64),
        .\CRC_OUT_reg[8]_0 (crcmodule_n_65),
        .\CRC_OUT_reg[8]_1 (crcmodule_n_74),
        .\CRC_OUT_reg[8]_2 (crcmodule_n_55),
        .\CRC_OUT_reg[9] (crcmodule_n_72),
        .\CRC_OUT_reg[9]_0 (crcmodule_n_68),
        .\CRC_OUT_reg[9]_1 (crcmodule_n_47),
        .D({rx_rs_n_2,rx_rs_n_3,rx_rs_n_4,rx_rs_n_5,rx_rs_n_6,rx_rs_n_7}),
        .E(terminator_location0),
        .\FSM_sequential_fifo_state_reg[0]_0 (fifo_state),
        .Q({start_lt,start_da}),
        .SS(datapath_main_n_80),
        .bad_frame_get(bad_frame_get),
        .bad_frame_get_reg(rx_bad_frame),
        .\bytes_cnt_reg[1] (bytes_cnt),
        .\bytes_cnt_reg[2] (crcmodule_n_4),
        .check_reset(check_reset),
        .check_reset_reg_0(statemachine_n_20),
        .clk_i(clk_i),
        .\da_addr_reg[40]_0 (datapath_main_n_195),
        .\da_addr_reg[6]_0 (datapath_main_n_194),
        .do_crc_check_reg(crcmodule_n_9),
        .\get_e_chk_reg[7]_0 (p_16_out),
        .get_error_code(get_error_code),
        .get_error_code_reg_0(statemachine_n_19),
        .get_sfd(get_sfd),
        .get_sfd0(get_sfd0),
        .get_terminator(get_terminator),
        .get_terminator_d1(get_terminator_d1),
        .get_terminator_d2(get_terminator_d2),
        .get_terminator_d2_reg(datapath_main_n_79),
        .get_terminator_d3(get_terminator_d3),
        .get_terminator_reg_0(datapath_main_n_73),
        .good_frame_get(good_frame_get),
        .good_frame_get_reg(rx_good_frame),
        .in0(in0[13]),
        .inband_fcs(inband_fcs),
        .qvDataOut({rxc8,rxd64}),
        .receiving(receiving),
        .recv_rst(recv_rst),
        .reset_dcm(reset_dcm),
        .rst_i(rst_i),
        .\rx_data_reg[63]_0 (rx_data),
        .\rx_data_valid_reg[7]_0 (rx_data_valid),
        .rxd64_d3(rxd64_d3),
        .\rxd64_d3_reg[20]_0 (datapath_main_n_113),
        .\rxd64_d3_reg[29]_0 (datapath_main_n_117),
        .\rxd64_d3_reg[30]_0 (datapath_main_n_112),
        .\rxd64_d3_reg[34]_0 (datapath_main_n_114),
        .\rxd64_d3_reg[40]_0 (datapath_main_n_120),
        .\rxd64_d3_reg[8]_0 (datapath_main_n_119),
        .\rxd64_d3_reg[9]_0 (datapath_main_n_121),
        .tagged_frame(tagged_frame),
        .tagged_frame_reg_0(rx_rs_n_95),
        .\terminator_location_reg[1]_0 ({datapath_main_n_74,datapath_main_n_75}),
        .\terminator_location_reg[2]_0 (terminator_location),
        .\terminator_location_reg[2]_1 ({rx_rs_n_83,rx_rs_n_84,rx_rs_n_85}),
        .this_cycle(this_cycle),
        .wait_crc_check(wait_crc_check));
  FDCE #(
    .INIT(1'b0)) 
    inband_fcs_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg_n_0_[50] ),
        .Q(inband_fcs));
  FDCE #(
    .INIT(1'b0)) 
    jumbo_enable_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg_n_0_[51] ),
        .Q(jumbo_enable));
  switch_elements_rxLenTypChecker lenchecker
       (.D({lenchecker_n_8,lenchecker_n_9}),
        .Q({statemachine_n_13,statemachine_n_14}),
        .bad_frame_get0(bad_frame_get0),
        .bad_frame_get_reg(crc_check_invalid),
        .clk_i(clk_i),
        .get_error_code(get_error_code),
        .get_terminator(get_terminator),
        .jumbo_enable(jumbo_enable),
        .jumbo_frame(jumbo_frame),
        .jumbo_frame0(jumbo_frame0),
        .large_error(large_error),
        .large_error_i_4(counters_n_12),
        .large_error_i_4_0(counters_n_14),
        .large_error_reg_0(counters_n_8),
        .large_error_reg_1(counters_n_11),
        .large_error_reg_2(counters_n_21),
        .length_128_255(length_128_255),
        .length_128_2550(length_128_2550),
        .length_256_511(length_256_511),
        .length_256_5110(length_256_5110),
        .length_512_1023(length_512_1023),
        .length_512_10230(length_512_10230),
        .length_65_127(length_65_127),
        .length_65_1270(length_65_1270),
        .\location_reg_reg[0]_0 (lenchecker_n_11),
        .\location_reg_reg[0]_1 (lenchecker_n_13),
        .\location_reg_reg[2]_0 (location_reg),
        .\location_reg_reg[2]_1 (terminator_location),
        .padded_frame(padded_frame),
        .padded_frame0(padded_frame0),
        .reset_dcm(reset_dcm),
        .small_error(small_error),
        .small_error0(small_error0),
        .tagged_frame(tagged_frame),
        .vlan_enable(vlan_enable));
  FDCE #(
    .INIT(1'b0)) 
    recv_enable_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg_n_0_[49] ),
        .Q(recv_enable));
  FDCE #(
    .INIT(1'b0)) 
    recv_rst_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg_n_0_[52] ),
        .Q(recv_rst));
  LUT2 #(
    .INIT(4'h1)) 
    rxCfgofRS_inferred_i_1
       (.I0(recv_rst),
        .I1(rst_i),
        .O(rxCfgofRS[2]));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT2 #(
    .INIT(4'h8)) 
    rxCfgofRS_inferred_i_2
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(rxCfgofRS[1]));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT2 #(
    .INIT(4'h2)) 
    rxCfgofRS_inferred_i_3
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(rxCfgofRS[0]));
  switch_elements_rxRSLayer rx_rs
       (.D({rx_rs_n_2,rx_rs_n_3,rx_rs_n_4,rx_rs_n_5,rx_rs_n_6,rx_rs_n_7}),
        .E(terminator_location0),
        .Q({rxc8,rxd64}),
        .clk_i(clk_i),
        .get_sfd0(get_sfd0),
        .\link_fault_reg[1] (Q),
        .\qvDataOut_reg[45] (rx_rs_n_95),
        .\qvDataOut_reg[62] (p_16_out),
        .\qvDataOut_reg[69] ({rx_rs_n_83,rx_rs_n_84,rx_rs_n_85}),
        .recv_rst(recv_rst),
        .reset_dcm(reset_dcm),
        .rst_i(rst_i),
        .\rxc4_in_tmp_reg[3] (\rxc4_in_tmp_reg[3] ),
        .rxclk_180(rxclk_180),
        .\rxd32_in_tmp_reg[31] (D),
        .this_cycle(this_cycle));
  switch_elements_rxStatModule rx_stat
       (.D({rxStatRegPlus_tmp09_out,small_error,rxStatRegPlus_tmp08_out,large_error,rxStatRegPlus_tmp05_out,rxStatRegPlus_tmp04_out,rxStatRegPlus_tmp03_out,rxStatRegPlus_tmp02_out,rxStatRegPlus_tmp01_out,rxStatRegPlus_tmp00_out,rxStatRegPlus_tmp0,crc_check_invalid,good_frame_get}),
        .clk_i(clk_i),
        .in0(in0[12:0]),
        .reset_dcm(reset_dcm));
  switch_elements_rxStateMachine statemachine
       (.D({rxStatRegPlus_tmp09_out,rxStatRegPlus_tmp08_out,rxStatRegPlus_tmp05_out,rxStatRegPlus_tmp04_out,rxStatRegPlus_tmp03_out,rxStatRegPlus_tmp02_out,rxStatRegPlus_tmp01_out,rxStatRegPlus_tmp00_out,rxStatRegPlus_tmp0,good_frame_get}),
        .\FSM_onehot_rxstate_reg[1]_0 (statemachine_n_19),
        .\FSM_onehot_rxstate_reg[3]_0 (statemachine_n_22),
        .\FSM_onehot_rxstate_reg[3]_1 (statemachine_n_23),
        .\FSM_onehot_rxstate_reg[3]_2 (statemachine_n_24),
        .\FSM_onehot_rxstate_reg[3]_3 (statemachine_n_25),
        .\FSM_onehot_rxstate_reg[5]_0 ({lenchecker_n_8,lenchecker_n_9}),
        .\FSM_sequential_fifo_state_reg[0] (statemachine_n_20),
        .Q({statemachine_n_13,statemachine_n_14,start_lt,start_da}),
        .bad_frame_get(bad_frame_get),
        .bad_frame_get0(bad_frame_get0),
        .bad_frame_get_reg_0({small_error,large_error}),
        .broad_valid(broad_valid),
        .check_reset(check_reset),
        .check_reset_reg(fifo_state),
        .clk_i(clk_i),
        .crc_64_en(crc_64_en),
        .do_crc_check(do_crc_check),
        .get_error_code(get_error_code),
        .get_sfd(get_sfd),
        .get_terminator(get_terminator),
        .good_frame_get_reg_0(crcmodule_n_5),
        .in0(in0[13]),
        .jumbo_frame(jumbo_frame),
        .length_128_255(length_128_255),
        .length_256_511(length_256_511),
        .length_512_1023(length_512_1023),
        .length_65_127(length_65_127),
        .multi_valid(multi_valid),
        .padded_frame(padded_frame),
        .receiving(receiving),
        .recv_enable(recv_enable),
        .reset_dcm(reset_dcm),
        .\value_reg[0] (statemachine_n_21),
        .\value_reg[10] ({frame_cnt[10],frame_cnt[7:4],frame_cnt[1:0]}),
        .\value_reg[10]_0 (counters_n_7),
        .\value_reg[1] (p_0_in),
        .\value_reg[5] (counters_n_13),
        .\value_reg[6] (counters_n_9),
        .wait_crc_check(wait_crc_check));
  FDCE #(
    .INIT(1'b0)) 
    vlan_enable_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\cfgRxRegData_reg_n_0_[48] ),
        .Q(vlan_enable));
endmodule

(* ORIG_REF_NAME = "rxStatModule" *) 
module switch_elements_rxStatModule
   (in0,
    D,
    clk_i,
    reset_dcm);
  output [12:0]in0;
  input [12:0]D;
  input clk_i;
  input reset_dcm;

  wire [12:0]D;
  wire clk_i;
  wire [12:0]in0;
  wire reset_dcm;

  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[0]),
        .Q(in0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[9]),
        .Q(in0[9]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[10]),
        .Q(in0[10]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[11]),
        .Q(in0[11]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[12]),
        .Q(in0[12]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[1]),
        .Q(in0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[2]),
        .Q(in0[2]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[3]),
        .Q(in0[3]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[4]),
        .Q(in0[4]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[5]),
        .Q(in0[5]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[6]),
        .Q(in0[6]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[7]),
        .Q(in0[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rxStatRegPlus_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(D[8]),
        .Q(in0[8]));
endmodule

(* ORIG_REF_NAME = "rxStateMachine" *) 
module switch_elements_rxStateMachine
   (D,
    bad_frame_get,
    wait_crc_check,
    crc_64_en,
    Q,
    \value_reg[1] ,
    receiving,
    \FSM_onehot_rxstate_reg[1]_0 ,
    \FSM_sequential_fifo_state_reg[0] ,
    \value_reg[0] ,
    \FSM_onehot_rxstate_reg[3]_0 ,
    \FSM_onehot_rxstate_reg[3]_1 ,
    \FSM_onehot_rxstate_reg[3]_2 ,
    \FSM_onehot_rxstate_reg[3]_3 ,
    good_frame_get_reg_0,
    clk_i,
    reset_dcm,
    bad_frame_get0,
    in0,
    get_error_code,
    \value_reg[10] ,
    get_terminator,
    bad_frame_get_reg_0,
    jumbo_frame,
    length_512_1023,
    length_256_511,
    length_128_255,
    length_65_127,
    padded_frame,
    multi_valid,
    broad_valid,
    check_reset_reg,
    get_sfd,
    recv_enable,
    \value_reg[5] ,
    \value_reg[6] ,
    \value_reg[10]_0 ,
    do_crc_check,
    check_reset,
    \FSM_onehot_rxstate_reg[5]_0 );
  output [9:0]D;
  output bad_frame_get;
  output wait_crc_check;
  output crc_64_en;
  output [3:0]Q;
  output [0:0]\value_reg[1] ;
  output receiving;
  output \FSM_onehot_rxstate_reg[1]_0 ;
  output \FSM_sequential_fifo_state_reg[0] ;
  output \value_reg[0] ;
  output \FSM_onehot_rxstate_reg[3]_0 ;
  output \FSM_onehot_rxstate_reg[3]_1 ;
  output \FSM_onehot_rxstate_reg[3]_2 ;
  output \FSM_onehot_rxstate_reg[3]_3 ;
  input good_frame_get_reg_0;
  input clk_i;
  input reset_dcm;
  input bad_frame_get0;
  input [0:0]in0;
  input get_error_code;
  input [6:0]\value_reg[10] ;
  input get_terminator;
  input [1:0]bad_frame_get_reg_0;
  input jumbo_frame;
  input length_512_1023;
  input length_256_511;
  input length_128_255;
  input length_65_127;
  input padded_frame;
  input multi_valid;
  input broad_valid;
  input [0:0]check_reset_reg;
  input get_sfd;
  input recv_enable;
  input \value_reg[5] ;
  input \value_reg[6] ;
  input \value_reg[10]_0 ;
  input do_crc_check;
  input check_reset;
  input [1:0]\FSM_onehot_rxstate_reg[5]_0 ;

  wire [9:0]D;
  wire \FSM_onehot_rxstate_next_reg[0]_i_1_n_0 ;
  wire \FSM_onehot_rxstate_next_reg[1]_i_1_n_0 ;
  wire \FSM_onehot_rxstate_next_reg[3]_i_1_n_0 ;
  wire \FSM_onehot_rxstate_next_reg_n_0_[0] ;
  wire \FSM_onehot_rxstate_next_reg_n_0_[1] ;
  wire \FSM_onehot_rxstate_next_reg_n_0_[2] ;
  wire \FSM_onehot_rxstate_next_reg_n_0_[3] ;
  wire \FSM_onehot_rxstate_next_reg_n_0_[4] ;
  wire \FSM_onehot_rxstate_next_reg_n_0_[5] ;
  wire \FSM_onehot_rxstate_reg[1]_0 ;
  wire \FSM_onehot_rxstate_reg[3]_0 ;
  wire \FSM_onehot_rxstate_reg[3]_1 ;
  wire \FSM_onehot_rxstate_reg[3]_2 ;
  wire \FSM_onehot_rxstate_reg[3]_3 ;
  wire [1:0]\FSM_onehot_rxstate_reg[5]_0 ;
  wire \FSM_onehot_rxstate_reg_n_0_[0] ;
  wire \FSM_sequential_fifo_state_reg[0] ;
  wire [3:0]Q;
  wire bad_frame_get;
  wire bad_frame_get0;
  wire [1:0]bad_frame_get_reg_0;
  wire broad_valid;
  wire check_reset;
  wire [0:0]check_reset_reg;
  wire clk_i;
  wire crc_64_en;
  wire do_crc_check;
  wire get_error_code;
  wire get_sfd;
  wire get_terminator;
  wire good_frame_get_i_1_n_0;
  wire good_frame_get_reg_0;
  wire [0:0]in0;
  wire jumbo_frame;
  wire length_128_255;
  wire length_256_511;
  wire length_512_1023;
  wire length_65_127;
  wire multi_valid;
  wire p_0_in;
  wire padded_frame;
  wire receiving;
  wire recv_enable;
  wire reset_dcm;
  wire rxstate_next;
  wire \value_reg[0] ;
  wire [6:0]\value_reg[10] ;
  wire \value_reg[10]_0 ;
  wire [0:0]\value_reg[1] ;
  wire \value_reg[5] ;
  wire \value_reg[6] ;
  wire wait_crc_check;
  wire wait_crc_check_i_1_n_0;

  (* XILINX_LEGACY_PRIM = "LDP" *) 
  LDPE #(
    .INIT(1'b1)) 
    \FSM_onehot_rxstate_next_reg[0] 
       (.D(\FSM_onehot_rxstate_next_reg[0]_i_1_n_0 ),
        .G(rxstate_next),
        .GE(1'b1),
        .PRE(reset_dcm),
        .Q(\FSM_onehot_rxstate_next_reg_n_0_[0] ));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT5 #(
    .INIT(32'h77777770)) 
    \FSM_onehot_rxstate_next_reg[0]_i_1 
       (.I0(get_sfd),
        .I1(recv_enable),
        .I2(p_0_in),
        .I3(Q[3]),
        .I4(\FSM_onehot_rxstate_reg_n_0_[0] ),
        .O(\FSM_onehot_rxstate_next_reg[0]_i_1_n_0 ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_next_reg[1] 
       (.CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg[1]_i_1_n_0 ),
        .G(rxstate_next),
        .GE(1'b1),
        .Q(\FSM_onehot_rxstate_next_reg_n_0_[1] ));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT5 #(
    .INIT(32'h88888880)) 
    \FSM_onehot_rxstate_next_reg[1]_i_1 
       (.I0(get_sfd),
        .I1(recv_enable),
        .I2(p_0_in),
        .I3(Q[3]),
        .I4(\FSM_onehot_rxstate_reg_n_0_[0] ),
        .O(\FSM_onehot_rxstate_next_reg[1]_i_1_n_0 ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_next_reg[2] 
       (.CLR(reset_dcm),
        .D(Q[0]),
        .G(rxstate_next),
        .GE(1'b1),
        .Q(\FSM_onehot_rxstate_next_reg_n_0_[2] ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_next_reg[3] 
       (.CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg[3]_i_1_n_0 ),
        .G(rxstate_next),
        .GE(1'b1),
        .Q(\FSM_onehot_rxstate_next_reg_n_0_[3] ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAABA)) 
    \FSM_onehot_rxstate_next_reg[3]_i_1 
       (.I0(Q[1]),
        .I1(get_terminator),
        .I2(Q[2]),
        .I3(get_error_code),
        .I4(bad_frame_get_reg_0[1]),
        .I5(bad_frame_get_reg_0[0]),
        .O(\FSM_onehot_rxstate_next_reg[3]_i_1_n_0 ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_next_reg[4] 
       (.CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_reg[5]_0 [0]),
        .G(rxstate_next),
        .GE(1'b1),
        .Q(\FSM_onehot_rxstate_next_reg_n_0_[4] ));
  (* XILINX_LEGACY_PRIM = "LDC" *) 
  LDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_next_reg[5] 
       (.CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_reg[5]_0 [1]),
        .G(rxstate_next),
        .GE(1'b1),
        .Q(\FSM_onehot_rxstate_next_reg_n_0_[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_onehot_rxstate_next_reg[5]_i_2 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(p_0_in),
        .I4(Q[3]),
        .I5(\FSM_onehot_rxstate_reg_n_0_[0] ),
        .O(rxstate_next));
  (* FSM_ENCODED_STATES = "rxReceiveLT:000100,rxGetError:010000,rxReceiveData:001000,rxIFGWait:100000,IDLE:000001,rxReceiveDA:000010" *) 
  FDPE #(
    .INIT(1'b1)) 
    \FSM_onehot_rxstate_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\FSM_onehot_rxstate_next_reg_n_0_[0] ),
        .PRE(reset_dcm),
        .Q(\FSM_onehot_rxstate_reg_n_0_[0] ));
  (* FSM_ENCODED_STATES = "rxReceiveLT:000100,rxGetError:010000,rxReceiveData:001000,rxIFGWait:100000,IDLE:000001,rxReceiveDA:000010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg_n_0_[1] ),
        .Q(Q[0]));
  (* FSM_ENCODED_STATES = "rxReceiveLT:000100,rxGetError:010000,rxReceiveData:001000,rxIFGWait:100000,IDLE:000001,rxReceiveDA:000010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg_n_0_[2] ),
        .Q(Q[1]));
  (* FSM_ENCODED_STATES = "rxReceiveLT:000100,rxGetError:010000,rxReceiveData:001000,rxIFGWait:100000,IDLE:000001,rxReceiveDA:000010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg_n_0_[3] ),
        .Q(Q[2]));
  (* FSM_ENCODED_STATES = "rxReceiveLT:000100,rxGetError:010000,rxReceiveData:001000,rxIFGWait:100000,IDLE:000001,rxReceiveDA:000010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg_n_0_[4] ),
        .Q(Q[3]));
  (* FSM_ENCODED_STATES = "rxReceiveLT:000100,rxGetError:010000,rxReceiveData:001000,rxIFGWait:100000,IDLE:000001,rxReceiveDA:000010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_onehot_rxstate_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(\FSM_onehot_rxstate_next_reg_n_0_[5] ),
        .Q(p_0_in));
  FDCE #(
    .INIT(1'b0)) 
    bad_frame_get_reg
       (.C(clk_i),
        .CE(good_frame_get_i_1_n_0),
        .CLR(reset_dcm),
        .D(bad_frame_get0),
        .Q(bad_frame_get));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'h54)) 
    check_reset_i_2
       (.I0(check_reset_reg),
        .I1(bad_frame_get),
        .I2(D[0]),
        .O(\FSM_sequential_fifo_state_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT5 #(
    .INIT(32'h0000AAA8)) 
    crc_64_en_i_1
       (.I0(in0),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(get_error_code),
        .O(crc_64_en));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'h01)) 
    get_error_code_i_2
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(\FSM_onehot_rxstate_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    good_frame_get_i_1
       (.I0(do_crc_check),
        .I1(wait_crc_check),
        .I2(bad_frame_get_reg_0[0]),
        .I3(bad_frame_get_reg_0[1]),
        .I4(check_reset),
        .I5(Q[3]),
        .O(good_frame_get_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    good_frame_get_reg
       (.C(clk_i),
        .CE(good_frame_get_i_1_n_0),
        .CLR(reset_dcm),
        .D(good_frame_get_reg_0),
        .Q(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    receiving_d1_i_1
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(receiving));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[14]_i_1 
       (.I0(D[0]),
        .I1(jumbo_frame),
        .O(D[8]));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT4 #(
    .INIT(16'hAAA8)) 
    \rxStatRegPlus[16]_i_1 
       (.I0(get_error_code),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(D[9]));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[2]_i_1 
       (.I0(D[0]),
        .I1(broad_valid),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[3]_i_1 
       (.I0(D[0]),
        .I1(multi_valid),
        .O(D[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[4]_i_1 
       (.I0(D[0]),
        .I1(padded_frame),
        .O(D[3]));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[5]_i_1 
       (.I0(D[0]),
        .I1(length_65_127),
        .O(D[4]));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[6]_i_1 
       (.I0(D[0]),
        .I1(length_128_255),
        .O(D[5]));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[7]_i_1 
       (.I0(D[0]),
        .I1(length_256_511),
        .O(D[6]));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rxStatRegPlus[8]_i_1 
       (.I0(D[0]),
        .I1(length_512_1023),
        .O(D[7]));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT4 #(
    .INIT(16'h5554)) 
    \value[0]_i_1 
       (.I0(\value_reg[10] [0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\value_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT5 #(
    .INIT(32'h00FEFE00)) 
    \value[10]_i_1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(\value_reg[10]_0 ),
        .I4(\value_reg[10] [6]),
        .O(\FSM_onehot_rxstate_reg[3]_3 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT5 #(
    .INIT(32'h66666660)) 
    \value[1]_i_1 
       (.I0(\value_reg[10] [1]),
        .I1(\value_reg[10] [0]),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(Q[0]),
        .O(\value_reg[1] ));
  LUT6 #(
    .INIT(64'hFE00FEFE00FE0000)) 
    \value[5]_i_1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(\value_reg[5] ),
        .I4(\value_reg[10] [2]),
        .I5(\value_reg[10] [3]),
        .O(\FSM_onehot_rxstate_reg[3]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT5 #(
    .INIT(32'hFE0000FE)) 
    \value[6]_i_1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(\value_reg[6] ),
        .I4(\value_reg[10] [4]),
        .O(\FSM_onehot_rxstate_reg[3]_1 ));
  LUT6 #(
    .INIT(64'hFE00FEFE00FE0000)) 
    \value[7]_i_1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(\value_reg[6] ),
        .I4(\value_reg[10] [4]),
        .I5(\value_reg[10] [5]),
        .O(\FSM_onehot_rxstate_reg[3]_2 ));
  LUT5 #(
    .INIT(32'hFFFF0004)) 
    wait_crc_check_i_1
       (.I0(do_crc_check),
        .I1(wait_crc_check),
        .I2(bad_frame_get_reg_0[0]),
        .I3(bad_frame_get_reg_0[1]),
        .I4(p_0_in),
        .O(wait_crc_check_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    wait_crc_check_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(reset_dcm),
        .D(wait_crc_check_i_1_n_0),
        .Q(wait_crc_check));
endmodule

(* ORIG_REF_NAME = "simple_spi_top" *) 
module switch_elements_simple_spi_top
   (ack_o,
    in0,
    sck_o,
    treg,
    dat_o,
    clk_i,
    E,
    out,
    \dat_o_reg[3]_0 ,
    dat_i,
    \treg_reg[0]_0 ,
    rst_i,
    \sper_reg[0]_0 ,
    \sper_reg[0]_1 );
  output ack_o;
  output in0;
  output sck_o;
  output [0:0]treg;
  output [7:0]dat_o;
  input clk_i;
  input [0:0]E;
  input out;
  input [1:0]\dat_o_reg[3]_0 ;
  input [7:0]dat_i;
  input \treg_reg[0]_0 ;
  input rst_i;
  input \sper_reg[0]_0 ;
  input \sper_reg[0]_1 ;

  wire [0:0]E;
  wire \FSM_sequential_state[0]_i_1_n_0 ;
  wire \FSM_sequential_state[1]_i_1_n_0 ;
  wire \FSM_sequential_state[1]_i_3_n_0 ;
  wire \FSM_sequential_state[1]_i_6_n_0 ;
  wire \FSM_sequential_state[1]_i_7_n_0 ;
  wire ack_o;
  wire ack_o0;
  wire [2:0]bcnt;
  wire \bcnt_reg_n_0_[0] ;
  wire \bcnt_reg_n_0_[1] ;
  wire \bcnt_reg_n_0_[2] ;
  wire clk_i;
  wire \clkcnt[11]_i_1_n_0 ;
  wire \clkcnt[11]_i_2_n_0 ;
  wire \clkcnt[11]_i_3_n_0 ;
  wire \clkcnt[2]_i_2_n_0 ;
  wire \clkcnt[3]_i_2_n_0 ;
  wire \clkcnt[4]_i_2_n_0 ;
  wire \clkcnt[5]_i_2_n_0 ;
  wire \clkcnt[6]_i_2_n_0 ;
  wire \clkcnt[7]_i_2_n_0 ;
  wire \clkcnt[8]_i_2_n_0 ;
  wire \clkcnt[9]_i_2_n_0 ;
  wire [11:0]clkcnt_reg;
  wire cpha;
  wire cpol;
  wire [7:0]dat_i;
  wire [7:0]dat_o;
  wire [1:0]\dat_o_reg[3]_0 ;
  wire [4:3]dout__0;
  wire [1:0]icnt;
  wire in0;
  wire inta_o0;
  wire out;
  wire p_0_in;
  wire [7:0]p_0_in__0;
  wire [10:0]p_0_in__1;
  wire p_7_in;
  wire rfifo_n_2;
  wire rfwe;
  wire rfwe_reg_n_0;
  wire rst_i;
  wire sck_o;
  wire sck_o_i_3_n_0;
  wire [3:0]sel0;
  wire spcr;
  wire \spcr_reg_n_0_[5] ;
  wire spe;
  wire sper;
  wire \sper_reg[0]_0 ;
  wire \sper_reg[0]_1 ;
  wire \sper_reg_n_0_[2] ;
  wire \sper_reg_n_0_[3] ;
  wire \sper_reg_n_0_[4] ;
  wire \sper_reg_n_0_[5] ;
  wire spie;
  wire spif;
  wire spif0;
  wire [1:0]state;
  wire [1:0]tcnt;
  wire \tcnt[0]_i_1_n_0 ;
  wire \tcnt[1]_i_1_n_0 ;
  wire [0:0]treg;
  wire [7:0]treg0_out;
  wire \treg[7]_i_1_n_0 ;
  wire [6:0]treg_0;
  wire \treg_reg[0]_0 ;
  wire wcol;
  wire wcol0;
  wire wfifo_n_0;
  wire wfifo_n_1;
  wire wfifo_n_13;
  wire wfre_reg_n_0;

  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'h55545555)) 
    \FSM_sequential_state[0]_i_1 
       (.I0(state[0]),
        .I1(\bcnt_reg_n_0_[0] ),
        .I2(\bcnt_reg_n_0_[2] ),
        .I3(\bcnt_reg_n_0_[1] ),
        .I4(state[1]),
        .O(\FSM_sequential_state[0]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_state[1]_i_1 
       (.I0(spe),
        .O(\FSM_sequential_state[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \FSM_sequential_state[1]_i_3 
       (.I0(state[1]),
        .I1(state[0]),
        .I2(p_0_in),
        .O(\FSM_sequential_state[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \FSM_sequential_state[1]_i_5 
       (.I0(clkcnt_reg[2]),
        .I1(clkcnt_reg[3]),
        .I2(clkcnt_reg[0]),
        .I3(clkcnt_reg[1]),
        .I4(\FSM_sequential_state[1]_i_6_n_0 ),
        .I5(\FSM_sequential_state[1]_i_7_n_0 ),
        .O(p_0_in));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \FSM_sequential_state[1]_i_6 
       (.I0(clkcnt_reg[9]),
        .I1(clkcnt_reg[8]),
        .I2(clkcnt_reg[11]),
        .I3(clkcnt_reg[10]),
        .O(\FSM_sequential_state[1]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \FSM_sequential_state[1]_i_7 
       (.I0(clkcnt_reg[5]),
        .I1(clkcnt_reg[4]),
        .I2(clkcnt_reg[7]),
        .I3(clkcnt_reg[6]),
        .O(\FSM_sequential_state[1]_i_7_n_0 ));
  (* FSM_ENCODED_STATES = "iSTATE:10,iSTATE0:10,iSTATE1:00,iSTATE2:01" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[0] 
       (.C(clk_i),
        .CE(wfifo_n_13),
        .D(\FSM_sequential_state[0]_i_1_n_0 ),
        .Q(state[0]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  (* FSM_ENCODED_STATES = "iSTATE:10,iSTATE0:10,iSTATE1:00,iSTATE2:01" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[1] 
       (.C(clk_i),
        .CE(wfifo_n_13),
        .D(\FSM_sequential_state[1]_i_3_n_0 ),
        .Q(state[1]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    ack_o_i_1
       (.I0(\sper_reg[0]_1 ),
        .I1(\sper_reg[0]_0 ),
        .I2(ack_o),
        .O(ack_o0));
  FDCE #(
    .INIT(1'b0)) 
    ack_o_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(E),
        .D(ack_o0),
        .Q(ack_o));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \bcnt[0]_i_1 
       (.I0(\bcnt_reg_n_0_[0] ),
        .I1(state[1]),
        .O(bcnt[0]));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT3 #(
    .INIT(8'h9F)) 
    \bcnt[1]_i_1 
       (.I0(\bcnt_reg_n_0_[0] ),
        .I1(\bcnt_reg_n_0_[1] ),
        .I2(state[1]),
        .O(bcnt[1]));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'hE1FF)) 
    \bcnt[2]_i_1 
       (.I0(\bcnt_reg_n_0_[1] ),
        .I1(\bcnt_reg_n_0_[0] ),
        .I2(\bcnt_reg_n_0_[2] ),
        .I3(state[1]),
        .O(bcnt[2]));
  FDRE #(
    .INIT(1'b0)) 
    \bcnt_reg[0] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(bcnt[0]),
        .Q(\bcnt_reg_n_0_[0] ),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \bcnt_reg[1] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(bcnt[1]),
        .Q(\bcnt_reg_n_0_[1] ),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \bcnt_reg[2] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(bcnt[2]),
        .Q(\bcnt_reg_n_0_[2] ),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFE0000FFFEFFFF)) 
    \clkcnt[0]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[1]),
        .I2(sel0[0]),
        .I3(sel0[2]),
        .I4(\clkcnt[11]_i_2_n_0 ),
        .I5(clkcnt_reg[0]),
        .O(p_0_in__1[0]));
  LUT6 #(
    .INIT(64'h80FF8000800080FF)) 
    \clkcnt[10]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[0]),
        .I2(sel0[1]),
        .I3(\clkcnt[11]_i_2_n_0 ),
        .I4(\clkcnt[11]_i_3_n_0 ),
        .I5(clkcnt_reg[10]),
        .O(p_0_in__1[10]));
  LUT4 #(
    .INIT(16'h4441)) 
    \clkcnt[11]_i_1 
       (.I0(\clkcnt[11]_i_2_n_0 ),
        .I1(clkcnt_reg[11]),
        .I2(\clkcnt[11]_i_3_n_0 ),
        .I3(clkcnt_reg[10]),
        .O(\clkcnt[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT4 #(
    .INIT(16'hFDDF)) 
    \clkcnt[11]_i_2 
       (.I0(spe),
        .I1(p_0_in),
        .I2(state[0]),
        .I3(state[1]),
        .O(\clkcnt[11]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \clkcnt[11]_i_3 
       (.I0(clkcnt_reg[8]),
        .I1(clkcnt_reg[6]),
        .I2(\clkcnt[7]_i_2_n_0 ),
        .I3(clkcnt_reg[7]),
        .I4(clkcnt_reg[9]),
        .O(\clkcnt[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFE00FE00FEFF)) 
    \clkcnt[1]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[1]),
        .I2(sel0[2]),
        .I3(\clkcnt[11]_i_2_n_0 ),
        .I4(clkcnt_reg[0]),
        .I5(clkcnt_reg[1]),
        .O(p_0_in__1[1]));
  LUT6 #(
    .INIT(64'hFEFFFE00FE00FEFF)) 
    \clkcnt[2]_i_1 
       (.I0(sel0[3]),
        .I1(\clkcnt[6]_i_2_n_0 ),
        .I2(sel0[2]),
        .I3(\clkcnt[11]_i_2_n_0 ),
        .I4(\clkcnt[2]_i_2_n_0 ),
        .I5(clkcnt_reg[2]),
        .O(p_0_in__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \clkcnt[2]_i_2 
       (.I0(clkcnt_reg[0]),
        .I1(clkcnt_reg[1]),
        .O(\clkcnt[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFBEAFFFFFBEA0000)) 
    \clkcnt[3]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[0]),
        .I2(sel0[1]),
        .I3(sel0[2]),
        .I4(\clkcnt[11]_i_2_n_0 ),
        .I5(\clkcnt[3]_i_2_n_0 ),
        .O(p_0_in__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT4 #(
    .INIT(16'hFE01)) 
    \clkcnt[3]_i_2 
       (.I0(clkcnt_reg[2]),
        .I1(clkcnt_reg[0]),
        .I2(clkcnt_reg[1]),
        .I3(clkcnt_reg[3]),
        .O(\clkcnt[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAFFFFEFAA0000)) 
    \clkcnt[4]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[1]),
        .I2(sel0[0]),
        .I3(sel0[2]),
        .I4(\clkcnt[11]_i_2_n_0 ),
        .I5(\clkcnt[4]_i_2_n_0 ),
        .O(p_0_in__1[4]));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT5 #(
    .INIT(32'hFFFE0001)) 
    \clkcnt[4]_i_2 
       (.I0(clkcnt_reg[3]),
        .I1(clkcnt_reg[1]),
        .I2(clkcnt_reg[0]),
        .I3(clkcnt_reg[2]),
        .I4(clkcnt_reg[4]),
        .O(\clkcnt[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEA00EA00EAFF)) 
    \clkcnt[5]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[1]),
        .I2(sel0[2]),
        .I3(\clkcnt[11]_i_2_n_0 ),
        .I4(\clkcnt[5]_i_2_n_0 ),
        .I5(clkcnt_reg[5]),
        .O(p_0_in__1[5]));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \clkcnt[5]_i_2 
       (.I0(clkcnt_reg[3]),
        .I1(clkcnt_reg[1]),
        .I2(clkcnt_reg[0]),
        .I3(clkcnt_reg[2]),
        .I4(clkcnt_reg[4]),
        .O(\clkcnt[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEA00EA00EAFF)) 
    \clkcnt[6]_i_1 
       (.I0(sel0[3]),
        .I1(\clkcnt[6]_i_2_n_0 ),
        .I2(sel0[2]),
        .I3(\clkcnt[11]_i_2_n_0 ),
        .I4(\clkcnt[7]_i_2_n_0 ),
        .I5(clkcnt_reg[6]),
        .O(p_0_in__1[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \clkcnt[6]_i_2 
       (.I0(sel0[1]),
        .I1(sel0[0]),
        .O(\clkcnt[6]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT5 #(
    .INIT(32'hBBB8888B)) 
    \clkcnt[7]_i_1 
       (.I0(sel0[3]),
        .I1(\clkcnt[11]_i_2_n_0 ),
        .I2(clkcnt_reg[6]),
        .I3(\clkcnt[7]_i_2_n_0 ),
        .I4(clkcnt_reg[7]),
        .O(p_0_in__1[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \clkcnt[7]_i_2 
       (.I0(clkcnt_reg[4]),
        .I1(clkcnt_reg[2]),
        .I2(clkcnt_reg[0]),
        .I3(clkcnt_reg[1]),
        .I4(clkcnt_reg[3]),
        .I5(clkcnt_reg[5]),
        .O(\clkcnt[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8FFA800A800A8FF)) 
    \clkcnt[8]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[0]),
        .I2(sel0[1]),
        .I3(\clkcnt[11]_i_2_n_0 ),
        .I4(\clkcnt[8]_i_2_n_0 ),
        .I5(clkcnt_reg[8]),
        .O(p_0_in__1[8]));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \clkcnt[8]_i_2 
       (.I0(clkcnt_reg[6]),
        .I1(\clkcnt[7]_i_2_n_0 ),
        .I2(clkcnt_reg[7]),
        .O(\clkcnt[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8F80808F)) 
    \clkcnt[9]_i_1 
       (.I0(sel0[3]),
        .I1(sel0[1]),
        .I2(\clkcnt[11]_i_2_n_0 ),
        .I3(\clkcnt[9]_i_2_n_0 ),
        .I4(clkcnt_reg[9]),
        .O(p_0_in__1[9]));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \clkcnt[9]_i_2 
       (.I0(clkcnt_reg[7]),
        .I1(\clkcnt[7]_i_2_n_0 ),
        .I2(clkcnt_reg[6]),
        .I3(clkcnt_reg[8]),
        .O(\clkcnt[9]_i_2_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[0]),
        .Q(clkcnt_reg[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[10]),
        .Q(clkcnt_reg[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\clkcnt[11]_i_1_n_0 ),
        .Q(clkcnt_reg[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[1]),
        .Q(clkcnt_reg[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[2]),
        .Q(clkcnt_reg[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[3]),
        .Q(clkcnt_reg[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[4]),
        .Q(clkcnt_reg[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[5]),
        .Q(clkcnt_reg[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[6]),
        .Q(clkcnt_reg[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[7]),
        .Q(clkcnt_reg[7]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[8]),
        .Q(clkcnt_reg[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \clkcnt_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__1[9]),
        .Q(clkcnt_reg[9]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[0]),
        .Q(dat_o[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[1]),
        .Q(dat_o[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[2]),
        .Q(dat_o[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[3]),
        .Q(dat_o[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[4]),
        .Q(dat_o[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[5]),
        .Q(dat_o[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[6]),
        .Q(dat_o[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \dat_o_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in__0[7]),
        .Q(dat_o[7]),
        .R(1'b0));
  LUT2 #(
    .INIT(4'h8)) 
    inta_o_i_1
       (.I0(spif),
        .I1(spie),
        .O(inta_o0));
  FDRE #(
    .INIT(1'b0)) 
    inta_o_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(inta_o0),
        .Q(in0),
        .R(1'b0));
  switch_elements_fifo4 rfifo
       (.D({p_0_in__0[7:4],p_0_in__0[1:0]}),
        .DOB(dout__0),
        .E(rfifo_n_2),
        .Q({spie,spe,\spcr_reg_n_0_[5] ,sel0[1:0]}),
        .clk_i(clk_i),
        .\dat_o_reg[7] ({icnt,\sper_reg_n_0_[5] ,\sper_reg_n_0_[4] ,sel0[3:2]}),
        .out(out),
        .\rp_reg[0]_0 (E),
        .\rp_reg[1]_0 (\dat_o_reg[3]_0 ),
        .\rp_reg[1]_1 (ack_o),
        .\rp_reg[1]_2 (\sper_reg[0]_0 ),
        .\rp_reg[1]_3 (\sper_reg[0]_1 ),
        .rst_i(rst_i),
        .spif(spif),
        .treg({treg,treg_0}),
        .wcol(wcol),
        .\wp_reg[0]_0 (rfwe_reg_n_0));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    rfwe_i_1
       (.I0(state[0]),
        .I1(p_0_in),
        .I2(\bcnt_reg_n_0_[1] ),
        .I3(\bcnt_reg_n_0_[2] ),
        .I4(\bcnt_reg_n_0_[0] ),
        .I5(state[1]),
        .O(rfwe));
  FDRE #(
    .INIT(1'b0)) 
    rfwe_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(rfwe),
        .Q(rfwe_reg_n_0),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0002FFFE)) 
    sck_o_i_3
       (.I0(cpol),
        .I1(\bcnt_reg_n_0_[0] ),
        .I2(\bcnt_reg_n_0_[2] ),
        .I3(\bcnt_reg_n_0_[1] ),
        .I4(sck_o),
        .O(sck_o_i_3_n_0));
  FDRE #(
    .INIT(1'b0)) 
    sck_o_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(wfifo_n_0),
        .Q(sck_o),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \spcr[7]_i_1 
       (.I0(out),
        .I1(\sper_reg[0]_0 ),
        .I2(\sper_reg[0]_1 ),
        .I3(\dat_o_reg[3]_0 [1]),
        .I4(\dat_o_reg[3]_0 [0]),
        .O(spcr));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[0] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[0]),
        .Q(sel0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[1] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[1]),
        .Q(sel0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[2] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[2]),
        .Q(cpha));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[3] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[3]),
        .Q(cpol));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[5] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[5]),
        .Q(\spcr_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[6] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[6]),
        .Q(spe));
  FDCE #(
    .INIT(1'b0)) 
    \spcr_reg[7] 
       (.C(clk_i),
        .CE(spcr),
        .CLR(E),
        .D(dat_i[7]),
        .Q(spie));
  LUT5 #(
    .INIT(32'h80000000)) 
    \sper[7]_i_1 
       (.I0(out),
        .I1(\sper_reg[0]_0 ),
        .I2(\sper_reg[0]_1 ),
        .I3(\dat_o_reg[3]_0 [1]),
        .I4(\dat_o_reg[3]_0 [0]),
        .O(sper));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[0] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[0]),
        .Q(sel0[2]));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[1] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[1]),
        .Q(sel0[3]));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[2] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[2]),
        .Q(\sper_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[3] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[3]),
        .Q(\sper_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[4] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[4]),
        .Q(\sper_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[5] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[5]),
        .Q(\sper_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[6] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[6]),
        .Q(icnt[0]));
  FDCE #(
    .INIT(1'b0)) 
    \sper_reg[7] 
       (.C(clk_i),
        .CE(sper),
        .CLR(E),
        .D(dat_i[7]),
        .Q(icnt[1]));
  LUT6 #(
    .INIT(64'h0000ABAAABAAABAA)) 
    spif_i_1
       (.I0(spif),
        .I1(tcnt[1]),
        .I2(tcnt[0]),
        .I3(rfwe_reg_n_0),
        .I4(dat_i[7]),
        .I5(p_7_in),
        .O(spif0));
  FDRE #(
    .INIT(1'b0)) 
    spif_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(spif0),
        .Q(spif),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT4 #(
    .INIT(16'h5F40)) 
    \tcnt[0]_i_1 
       (.I0(tcnt[0]),
        .I1(tcnt[1]),
        .I2(spe),
        .I3(icnt[0]),
        .O(\tcnt[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT4 #(
    .INIT(16'h9F80)) 
    \tcnt[1]_i_1 
       (.I0(tcnt[0]),
        .I1(tcnt[1]),
        .I2(spe),
        .I3(icnt[1]),
        .O(\tcnt[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \tcnt_reg[0] 
       (.C(clk_i),
        .CE(rfifo_n_2),
        .D(\tcnt[0]_i_1_n_0 ),
        .Q(tcnt[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \tcnt_reg[1] 
       (.C(clk_i),
        .CE(rfifo_n_2),
        .D(\tcnt[1]_i_1_n_0 ),
        .Q(tcnt[1]),
        .R(1'b0));
  LUT3 #(
    .INIT(8'h45)) 
    \treg[7]_i_1 
       (.I0(state[0]),
        .I1(p_0_in),
        .I2(state[1]),
        .O(\treg[7]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[0] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[0]),
        .Q(treg_0[0]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[1] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[1]),
        .Q(treg_0[1]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[2] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[2]),
        .Q(treg_0[2]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[3] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[3]),
        .Q(treg_0[3]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[4] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[4]),
        .Q(treg_0[4]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[5] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[5]),
        .Q(treg_0[5]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[6] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[6]),
        .Q(treg_0[6]),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \treg_reg[7] 
       (.C(clk_i),
        .CE(\treg[7]_i_1_n_0 ),
        .D(treg0_out[7]),
        .Q(treg),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    wcol_i_3
       (.I0(out),
        .I1(\sper_reg[0]_0 ),
        .I2(\sper_reg[0]_1 ),
        .I3(\dat_o_reg[3]_0 [1]),
        .I4(\dat_o_reg[3]_0 [0]),
        .O(p_7_in));
  FDRE #(
    .INIT(1'b0)) 
    wcol_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(wcol0),
        .Q(wcol),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
  switch_elements_fifo4_5 wfifo
       (.D(treg0_out),
        .DOB(dout__0),
        .E(wfifo_n_13),
        .\FSM_sequential_state_reg[0] (wfifo_n_1),
        .\FSM_sequential_state_reg[1] (wfifo_n_0),
        .Q(state),
        .clk_i(clk_i),
        .dat_i(dat_i),
        .\dat_o_reg[3] ({\sper_reg_n_0_[3] ,\sper_reg_n_0_[2] }),
        .\dat_o_reg[3]_0 (\dat_o_reg[3]_0 ),
        .gb_reg_0({spe,cpol,cpha}),
        .gb_reg_1(wfre_reg_n_0),
        .out(out),
        .p_0_in(p_0_in),
        .p_7_in(p_7_in),
        .rst_i(rst_i),
        .sck_o_reg(sck_o_i_3_n_0),
        .sck_o_reg_0(sck_o),
        .\sper_reg[3] (p_0_in__0[3:2]),
        .\treg_reg[0] (\treg_reg[0]_0 ),
        .\treg_reg[7] (treg_0),
        .wcol(wcol),
        .wcol0(wcol0),
        .\wp_reg[0]_0 (E),
        .\wp_reg[1]_0 (ack_o),
        .\wp_reg[1]_1 (\sper_reg[0]_0 ),
        .\wp_reg[1]_2 (\sper_reg[0]_1 ));
  FDRE #(
    .INIT(1'b0)) 
    wfre_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(wfifo_n_1),
        .Q(wfre_reg_n_0),
        .R(\FSM_sequential_state[1]_i_1_n_0 ));
endmodule

(* ORIG_REF_NAME = "singleDouble" *) 
module switch_elements_singleDouble
   (CO,
    \count_zeros_reg[16]_0 ,
    \count_zeros_reg[16]_1 ,
    md16_nd,
    D,
    rst_i_0,
    rst_i_1,
    rst_i_2,
    in0,
    ce_i_d_reg_0,
    clk_i,
    rst_i,
    out,
    \FSM_sequential_state_reg[1] ,
    \FSM_sequential_state_reg[1]_0 ,
    Q,
    \FSM_sequential_state_reg[1]_1 ,
    \FSM_sequential_state_reg[1]_2 );
  output [0:0]CO;
  output [0:0]\count_zeros_reg[16]_0 ;
  output [0:0]\count_zeros_reg[16]_1 ;
  output md16_nd;
  output [0:0]D;
  output rst_i_0;
  output rst_i_1;
  output rst_i_2;
  output [3:0]in0;
  input ce_i_d_reg_0;
  input clk_i;
  input rst_i;
  input out;
  input \FSM_sequential_state_reg[1] ;
  input \FSM_sequential_state_reg[1]_0 ;
  input [0:0]Q;
  input \FSM_sequential_state_reg[1]_1 ;
  input \FSM_sequential_state_reg[1]_2 ;

  wire [0:0]CO;
  wire [0:0]D;
  wire \FSM_sequential_state[1]_i_2__0_n_0 ;
  wire \FSM_sequential_state[1]_i_3__0_n_0 ;
  wire \FSM_sequential_state[1]_i_4__0_n_0 ;
  wire \FSM_sequential_state_reg[1] ;
  wire \FSM_sequential_state_reg[1]_0 ;
  wire \FSM_sequential_state_reg[1]_1 ;
  wire \FSM_sequential_state_reg[1]_2 ;
  wire [0:0]Q;
  wire ce_i_d;
  wire ce_i_d2;
  wire ce_i_d_reg_0;
  wire clk_i;
  wire count_ones;
  wire \count_ones[0]_i_10_n_0 ;
  wire \count_ones[0]_i_11_n_0 ;
  wire \count_ones[0]_i_3_n_0 ;
  wire \count_ones[0]_i_4_n_0 ;
  wire \count_ones[0]_i_5_n_0 ;
  wire \count_ones[0]_i_6_n_0 ;
  wire \count_ones[0]_i_7_n_0 ;
  wire \count_ones[0]_i_8_n_0 ;
  wire \count_ones[0]_i_9_n_0 ;
  wire \count_ones[16]_i_2_n_0 ;
  wire \count_ones[8]_i_2_n_0 ;
  wire \count_ones[8]_i_3_n_0 ;
  wire \count_ones[8]_i_4_n_0 ;
  wire \count_ones[8]_i_5_n_0 ;
  wire \count_ones[8]_i_6_n_0 ;
  wire \count_ones[8]_i_7_n_0 ;
  wire \count_ones[8]_i_8_n_0 ;
  wire \count_ones[8]_i_9_n_0 ;
  wire [16:0]count_ones_reg;
  wire \count_ones_reg[0]_i_2_n_0 ;
  wire \count_ones_reg[0]_i_2_n_1 ;
  wire \count_ones_reg[0]_i_2_n_10 ;
  wire \count_ones_reg[0]_i_2_n_11 ;
  wire \count_ones_reg[0]_i_2_n_12 ;
  wire \count_ones_reg[0]_i_2_n_13 ;
  wire \count_ones_reg[0]_i_2_n_14 ;
  wire \count_ones_reg[0]_i_2_n_15 ;
  wire \count_ones_reg[0]_i_2_n_2 ;
  wire \count_ones_reg[0]_i_2_n_3 ;
  wire \count_ones_reg[0]_i_2_n_4 ;
  wire \count_ones_reg[0]_i_2_n_5 ;
  wire \count_ones_reg[0]_i_2_n_6 ;
  wire \count_ones_reg[0]_i_2_n_7 ;
  wire \count_ones_reg[0]_i_2_n_8 ;
  wire \count_ones_reg[0]_i_2_n_9 ;
  wire \count_ones_reg[16]_i_1_n_15 ;
  wire \count_ones_reg[8]_i_1_n_0 ;
  wire \count_ones_reg[8]_i_1_n_1 ;
  wire \count_ones_reg[8]_i_1_n_10 ;
  wire \count_ones_reg[8]_i_1_n_11 ;
  wire \count_ones_reg[8]_i_1_n_12 ;
  wire \count_ones_reg[8]_i_1_n_13 ;
  wire \count_ones_reg[8]_i_1_n_14 ;
  wire \count_ones_reg[8]_i_1_n_15 ;
  wire \count_ones_reg[8]_i_1_n_2 ;
  wire \count_ones_reg[8]_i_1_n_3 ;
  wire \count_ones_reg[8]_i_1_n_4 ;
  wire \count_ones_reg[8]_i_1_n_5 ;
  wire \count_ones_reg[8]_i_1_n_6 ;
  wire \count_ones_reg[8]_i_1_n_7 ;
  wire \count_ones_reg[8]_i_1_n_8 ;
  wire \count_ones_reg[8]_i_1_n_9 ;
  wire \count_zeros[0]_i_10_n_0 ;
  wire \count_zeros[0]_i_2_n_0 ;
  wire \count_zeros[0]_i_3_n_0 ;
  wire \count_zeros[0]_i_4_n_0 ;
  wire \count_zeros[0]_i_5_n_0 ;
  wire \count_zeros[0]_i_6_n_0 ;
  wire \count_zeros[0]_i_7_n_0 ;
  wire \count_zeros[0]_i_8_n_0 ;
  wire \count_zeros[0]_i_9_n_0 ;
  wire \count_zeros[16]_i_2_n_0 ;
  wire \count_zeros[8]_i_2_n_0 ;
  wire \count_zeros[8]_i_3_n_0 ;
  wire \count_zeros[8]_i_4_n_0 ;
  wire \count_zeros[8]_i_5_n_0 ;
  wire \count_zeros[8]_i_6_n_0 ;
  wire \count_zeros[8]_i_7_n_0 ;
  wire \count_zeros[8]_i_8_n_0 ;
  wire \count_zeros[8]_i_9_n_0 ;
  wire [16:0]count_zeros_reg;
  wire \count_zeros_reg[0]_i_1_n_0 ;
  wire \count_zeros_reg[0]_i_1_n_1 ;
  wire \count_zeros_reg[0]_i_1_n_10 ;
  wire \count_zeros_reg[0]_i_1_n_11 ;
  wire \count_zeros_reg[0]_i_1_n_12 ;
  wire \count_zeros_reg[0]_i_1_n_13 ;
  wire \count_zeros_reg[0]_i_1_n_14 ;
  wire \count_zeros_reg[0]_i_1_n_15 ;
  wire \count_zeros_reg[0]_i_1_n_2 ;
  wire \count_zeros_reg[0]_i_1_n_3 ;
  wire \count_zeros_reg[0]_i_1_n_4 ;
  wire \count_zeros_reg[0]_i_1_n_5 ;
  wire \count_zeros_reg[0]_i_1_n_6 ;
  wire \count_zeros_reg[0]_i_1_n_7 ;
  wire \count_zeros_reg[0]_i_1_n_8 ;
  wire \count_zeros_reg[0]_i_1_n_9 ;
  wire [0:0]\count_zeros_reg[16]_0 ;
  wire [0:0]\count_zeros_reg[16]_1 ;
  wire \count_zeros_reg[16]_i_1_n_15 ;
  wire \count_zeros_reg[8]_i_1_n_0 ;
  wire \count_zeros_reg[8]_i_1_n_1 ;
  wire \count_zeros_reg[8]_i_1_n_10 ;
  wire \count_zeros_reg[8]_i_1_n_11 ;
  wire \count_zeros_reg[8]_i_1_n_12 ;
  wire \count_zeros_reg[8]_i_1_n_13 ;
  wire \count_zeros_reg[8]_i_1_n_14 ;
  wire \count_zeros_reg[8]_i_1_n_15 ;
  wire \count_zeros_reg[8]_i_1_n_2 ;
  wire \count_zeros_reg[8]_i_1_n_3 ;
  wire \count_zeros_reg[8]_i_1_n_4 ;
  wire \count_zeros_reg[8]_i_1_n_5 ;
  wire \count_zeros_reg[8]_i_1_n_6 ;
  wire \count_zeros_reg[8]_i_1_n_7 ;
  wire \count_zeros_reg[8]_i_1_n_8 ;
  wire \count_zeros_reg[8]_i_1_n_9 ;
  wire [2:0]ct_state;
  wire \ct_state[1]_i_2_n_0 ;
  wire \ct_state[2]_i_3_n_0 ;
  wire \ct_state[2]_i_4_n_0 ;
  wire data_i_d;
  wire data_i_d2;
  wire double_one;
  wire i__carry__0_i_1__0_n_0;
  wire i__carry__0_i_1__1_n_0;
  wire i__carry__0_i_1_n_0;
  wire i__carry_i_10__0_n_0;
  wire i__carry_i_10__1_n_0;
  wire i__carry_i_10__4_n_0;
  wire i__carry_i_10_n_0;
  wire i__carry_i_11__0_n_0;
  wire i__carry_i_11__1_n_0;
  wire i__carry_i_11__2_n_0;
  wire i__carry_i_11__3_n_0;
  wire i__carry_i_12__1_n_0;
  wire i__carry_i_12__2_n_0;
  wire i__carry_i_12__3_n_0;
  wire i__carry_i_12_n_0;
  wire i__carry_i_13__0_n_0;
  wire i__carry_i_13__1_n_0;
  wire i__carry_i_13__2_n_0;
  wire i__carry_i_13__3_n_0;
  wire i__carry_i_14__0_n_0;
  wire i__carry_i_14__1_n_0;
  wire i__carry_i_15__0_n_0;
  wire i__carry_i_15__1_n_0;
  wire i__carry_i_1__0_n_0;
  wire i__carry_i_1__1_n_0;
  wire i__carry_i_1__4_n_0;
  wire i__carry_i_1_n_0;
  wire i__carry_i_2__0_n_0;
  wire i__carry_i_2__1_n_0;
  wire i__carry_i_2__4_n_0;
  wire i__carry_i_2_n_0;
  wire i__carry_i_3__0_n_0;
  wire i__carry_i_3__1_n_0;
  wire i__carry_i_3__4_n_0;
  wire i__carry_i_3_n_0;
  wire i__carry_i_4__0_n_0;
  wire i__carry_i_4__1_n_0;
  wire i__carry_i_4__4_n_0;
  wire i__carry_i_4_n_0;
  wire i__carry_i_5__0_n_0;
  wire i__carry_i_5__1_n_0;
  wire i__carry_i_5__4_n_0;
  wire i__carry_i_5_n_0;
  wire i__carry_i_6__0_n_0;
  wire i__carry_i_6__3_n_0;
  wire i__carry_i_6__4_n_0;
  wire i__carry_i_6_n_0;
  wire i__carry_i_7__0_n_0;
  wire i__carry_i_7__3_n_0;
  wire i__carry_i_7__4_n_0;
  wire i__carry_i_7_n_0;
  wire i__carry_i_8__2_n_0;
  wire i__carry_i_8__3_n_0;
  wire i__carry_i_8__4_n_0;
  wire i__carry_i_8_n_0;
  wire i__carry_i_9__0_n_0;
  wire i__carry_i_9__3_n_0;
  wire i__carry_i_9__4_n_0;
  wire i__carry_i_9_n_0;
  wire [3:0]in0;
  wire load;
  wire md16_nd;
  wire [2:0]nxt_state;
  wire out;
  wire q_o0_carry_i_10_n_0;
  wire q_o0_carry_i_11_n_0;
  wire q_o0_carry_i_12_n_0;
  wire q_o0_carry_i_13_n_0;
  wire q_o0_carry_i_14_n_0;
  wire q_o0_carry_i_15_n_0;
  wire q_o0_carry_i_1_n_0;
  wire q_o0_carry_i_2_n_0;
  wire q_o0_carry_i_3_n_0;
  wire q_o0_carry_i_4_n_0;
  wire q_o0_carry_i_5_n_0;
  wire q_o0_carry_i_6_n_0;
  wire q_o0_carry_i_7_n_0;
  wire q_o0_carry_i_8_n_0;
  wire q_o0_carry_i_9_n_0;
  wire q_o0_carry_n_0;
  wire q_o0_carry_n_1;
  wire q_o0_carry_n_2;
  wire q_o0_carry_n_3;
  wire q_o0_carry_n_4;
  wire q_o0_carry_n_5;
  wire q_o0_carry_n_6;
  wire q_o0_carry_n_7;
  wire \q_o0_inferred__0/i__carry_n_0 ;
  wire \q_o0_inferred__0/i__carry_n_1 ;
  wire \q_o0_inferred__0/i__carry_n_2 ;
  wire \q_o0_inferred__0/i__carry_n_3 ;
  wire \q_o0_inferred__0/i__carry_n_4 ;
  wire \q_o0_inferred__0/i__carry_n_5 ;
  wire \q_o0_inferred__0/i__carry_n_6 ;
  wire \q_o0_inferred__0/i__carry_n_7 ;
  wire q_o1;
  wire q_o10_in;
  wire q_o1_carry__0_i_1_n_0;
  wire q_o1_carry_i_10_n_0;
  wire q_o1_carry_i_11_n_0;
  wire q_o1_carry_i_12_n_0;
  wire q_o1_carry_i_13_n_0;
  wire q_o1_carry_i_14_n_0;
  wire q_o1_carry_i_15_n_0;
  wire q_o1_carry_i_1_n_0;
  wire q_o1_carry_i_2_n_0;
  wire q_o1_carry_i_3_n_0;
  wire q_o1_carry_i_4_n_0;
  wire q_o1_carry_i_5_n_0;
  wire q_o1_carry_i_6_n_0;
  wire q_o1_carry_i_7_n_0;
  wire q_o1_carry_i_8_n_0;
  wire q_o1_carry_i_9_n_0;
  wire q_o1_carry_n_0;
  wire q_o1_carry_n_1;
  wire q_o1_carry_n_2;
  wire q_o1_carry_n_3;
  wire q_o1_carry_n_4;
  wire q_o1_carry_n_5;
  wire q_o1_carry_n_6;
  wire q_o1_carry_n_7;
  wire \q_o1_inferred__0/i__carry_n_0 ;
  wire \q_o1_inferred__0/i__carry_n_1 ;
  wire \q_o1_inferred__0/i__carry_n_2 ;
  wire \q_o1_inferred__0/i__carry_n_3 ;
  wire \q_o1_inferred__0/i__carry_n_4 ;
  wire \q_o1_inferred__0/i__carry_n_5 ;
  wire \q_o1_inferred__0/i__carry_n_6 ;
  wire \q_o1_inferred__0/i__carry_n_7 ;
  wire \q_o1_inferred__1/i__carry_n_0 ;
  wire \q_o1_inferred__1/i__carry_n_1 ;
  wire \q_o1_inferred__1/i__carry_n_2 ;
  wire \q_o1_inferred__1/i__carry_n_3 ;
  wire \q_o1_inferred__1/i__carry_n_4 ;
  wire \q_o1_inferred__1/i__carry_n_5 ;
  wire \q_o1_inferred__1/i__carry_n_6 ;
  wire \q_o1_inferred__1/i__carry_n_7 ;
  wire \q_o1_inferred__2/i__carry_n_0 ;
  wire \q_o1_inferred__2/i__carry_n_1 ;
  wire \q_o1_inferred__2/i__carry_n_2 ;
  wire \q_o1_inferred__2/i__carry_n_3 ;
  wire \q_o1_inferred__2/i__carry_n_4 ;
  wire \q_o1_inferred__2/i__carry_n_5 ;
  wire \q_o1_inferred__2/i__carry_n_6 ;
  wire \q_o1_inferred__2/i__carry_n_7 ;
  wire rst_i;
  wire rst_i_0;
  wire rst_i_1;
  wire rst_i_2;
  wire [7:0]\NLW_count_ones_reg[16]_i_1_CO_UNCONNECTED ;
  wire [7:1]\NLW_count_ones_reg[16]_i_1_O_UNCONNECTED ;
  wire [7:0]\NLW_count_zeros_reg[16]_i_1_CO_UNCONNECTED ;
  wire [7:1]\NLW_count_zeros_reg[16]_i_1_O_UNCONNECTED ;
  wire [7:0]NLW_q_o0_carry_O_UNCONNECTED;
  wire [7:1]NLW_q_o0_carry__0_CO_UNCONNECTED;
  wire [7:0]NLW_q_o0_carry__0_O_UNCONNECTED;
  wire [7:0]\NLW_q_o0_inferred__0/i__carry_O_UNCONNECTED ;
  wire [7:1]\NLW_q_o0_inferred__0/i__carry__0_CO_UNCONNECTED ;
  wire [7:0]\NLW_q_o0_inferred__0/i__carry__0_O_UNCONNECTED ;
  wire [7:0]NLW_q_o1_carry_O_UNCONNECTED;
  wire [7:1]NLW_q_o1_carry__0_CO_UNCONNECTED;
  wire [7:0]NLW_q_o1_carry__0_O_UNCONNECTED;
  wire [7:0]\NLW_q_o1_inferred__0/i__carry_O_UNCONNECTED ;
  wire [7:1]\NLW_q_o1_inferred__0/i__carry__0_CO_UNCONNECTED ;
  wire [7:0]\NLW_q_o1_inferred__0/i__carry__0_O_UNCONNECTED ;
  wire [7:0]\NLW_q_o1_inferred__1/i__carry_O_UNCONNECTED ;
  wire [7:1]\NLW_q_o1_inferred__1/i__carry__0_CO_UNCONNECTED ;
  wire [7:0]\NLW_q_o1_inferred__1/i__carry__0_O_UNCONNECTED ;
  wire [7:0]\NLW_q_o1_inferred__2/i__carry_O_UNCONNECTED ;
  wire [7:1]\NLW_q_o1_inferred__2/i__carry__0_CO_UNCONNECTED ;
  wire [7:0]\NLW_q_o1_inferred__2/i__carry__0_O_UNCONNECTED ;

  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT4 #(
    .INIT(16'h0111)) 
    \FSM_sequential_state[0]_i_3 
       (.I0(rst_i),
        .I1(double_one),
        .I2(q_o1),
        .I3(q_o10_in),
        .O(rst_i_2));
  LUT6 #(
    .INIT(64'hFF00E000E000E000)) 
    \FSM_sequential_state[1]_i_1__0 
       (.I0(\FSM_sequential_state[1]_i_2__0_n_0 ),
        .I1(\FSM_sequential_state[1]_i_3__0_n_0 ),
        .I2(\FSM_sequential_state[1]_i_4__0_n_0 ),
        .I3(\FSM_sequential_state_reg[1] ),
        .I4(\FSM_sequential_state_reg[1]_0 ),
        .I5(Q),
        .O(D));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \FSM_sequential_state[1]_i_2__0 
       (.I0(double_one),
        .I1(rst_i),
        .I2(\FSM_sequential_state_reg[1]_1 ),
        .I3(\count_zeros_reg[16]_1 ),
        .I4(q_o10_in),
        .I5(q_o1),
        .O(\FSM_sequential_state[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0002020200000000)) 
    \FSM_sequential_state[1]_i_3__0 
       (.I0(\count_zeros_reg[16]_1 ),
        .I1(rst_i),
        .I2(double_one),
        .I3(q_o1),
        .I4(q_o10_in),
        .I5(\FSM_sequential_state_reg[1]_2 ),
        .O(\FSM_sequential_state[1]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \FSM_sequential_state[1]_i_4__0 
       (.I0(\count_zeros_reg[16]_0 ),
        .I1(CO),
        .O(\FSM_sequential_state[1]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'h4FF44444)) 
    \FSM_sequential_state[2]_i_2 
       (.I0(ce_i_d2),
        .I1(ce_i_d),
        .I2(data_i_d),
        .I3(data_i_d2),
        .I4(ce_i_d_reg_0),
        .O(md16_nd));
  LUT6 #(
    .INIT(64'h0007000000000000)) 
    \FSM_sequential_state[2]_i_4 
       (.I0(q_o10_in),
        .I1(q_o1),
        .I2(double_one),
        .I3(rst_i),
        .I4(CO),
        .I5(\count_zeros_reg[16]_0 ),
        .O(rst_i_1));
  LUT6 #(
    .INIT(64'h0000007000700070)) 
    \FSM_sequential_state[2]_i_5 
       (.I0(q_o10_in),
        .I1(q_o1),
        .I2(double_one),
        .I3(rst_i),
        .I4(CO),
        .I5(\count_zeros_reg[16]_0 ),
        .O(rst_i_0));
  FDCE #(
    .INIT(1'b0)) 
    ce_i_d2_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(ce_i_d),
        .Q(ce_i_d2));
  FDCE #(
    .INIT(1'b0)) 
    ce_i_d_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(ce_i_d_reg_0),
        .Q(ce_i_d));
  LUT3 #(
    .INIT(8'h12)) 
    \count_ones[0]_i_1 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .O(count_ones));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_10 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[1]),
        .O(\count_ones[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h5551)) 
    \count_ones[0]_i_11 
       (.I0(count_ones_reg[0]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_ones[0]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \count_ones[0]_i_3 
       (.I0(ct_state[2]),
        .I1(ct_state[0]),
        .I2(ct_state[1]),
        .O(\count_ones[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_4 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[7]),
        .O(\count_ones[0]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_5 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[6]),
        .O(\count_ones[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_6 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[5]),
        .O(\count_ones[0]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_7 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[4]),
        .O(\count_ones[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_8 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[3]),
        .O(\count_ones[0]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[0]_i_9 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[2]),
        .O(\count_ones[0]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[16]_i_2 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[16]),
        .O(\count_ones[16]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_2 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[15]),
        .O(\count_ones[8]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_3 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[14]),
        .O(\count_ones[8]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_4 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[13]),
        .O(\count_ones[8]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_5 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[12]),
        .O(\count_ones[8]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_6 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[11]),
        .O(\count_ones[8]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_7 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[10]),
        .O(\count_ones[8]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_8 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[9]),
        .O(\count_ones[8]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hFD00)) 
    \count_ones[8]_i_9 
       (.I0(ct_state[1]),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(count_ones_reg[8]),
        .O(\count_ones[8]_i_9_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[0] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_15 ),
        .Q(count_ones_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \count_ones_reg[0]_i_2 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\count_ones_reg[0]_i_2_n_0 ,\count_ones_reg[0]_i_2_n_1 ,\count_ones_reg[0]_i_2_n_2 ,\count_ones_reg[0]_i_2_n_3 ,\count_ones_reg[0]_i_2_n_4 ,\count_ones_reg[0]_i_2_n_5 ,\count_ones_reg[0]_i_2_n_6 ,\count_ones_reg[0]_i_2_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\count_ones[0]_i_3_n_0 }),
        .O({\count_ones_reg[0]_i_2_n_8 ,\count_ones_reg[0]_i_2_n_9 ,\count_ones_reg[0]_i_2_n_10 ,\count_ones_reg[0]_i_2_n_11 ,\count_ones_reg[0]_i_2_n_12 ,\count_ones_reg[0]_i_2_n_13 ,\count_ones_reg[0]_i_2_n_14 ,\count_ones_reg[0]_i_2_n_15 }),
        .S({\count_ones[0]_i_4_n_0 ,\count_ones[0]_i_5_n_0 ,\count_ones[0]_i_6_n_0 ,\count_ones[0]_i_7_n_0 ,\count_ones[0]_i_8_n_0 ,\count_ones[0]_i_9_n_0 ,\count_ones[0]_i_10_n_0 ,\count_ones[0]_i_11_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[10] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_13 ),
        .Q(count_ones_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[11] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_12 ),
        .Q(count_ones_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[12] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_11 ),
        .Q(count_ones_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[13] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_10 ),
        .Q(count_ones_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[14] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_9 ),
        .Q(count_ones_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[15] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_8 ),
        .Q(count_ones_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[16] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[16]_i_1_n_15 ),
        .Q(count_ones_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \count_ones_reg[16]_i_1 
       (.CI(\count_ones_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO(\NLW_count_ones_reg[16]_i_1_CO_UNCONNECTED [7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_count_ones_reg[16]_i_1_O_UNCONNECTED [7:1],\count_ones_reg[16]_i_1_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\count_ones[16]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[1] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_14 ),
        .Q(count_ones_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[2] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_13 ),
        .Q(count_ones_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[3] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_12 ),
        .Q(count_ones_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[4] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_11 ),
        .Q(count_ones_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[5] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_10 ),
        .Q(count_ones_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[6] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_9 ),
        .Q(count_ones_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[7] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[0]_i_2_n_8 ),
        .Q(count_ones_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[8] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_15 ),
        .Q(count_ones_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \count_ones_reg[8]_i_1 
       (.CI(\count_ones_reg[0]_i_2_n_0 ),
        .CI_TOP(1'b0),
        .CO({\count_ones_reg[8]_i_1_n_0 ,\count_ones_reg[8]_i_1_n_1 ,\count_ones_reg[8]_i_1_n_2 ,\count_ones_reg[8]_i_1_n_3 ,\count_ones_reg[8]_i_1_n_4 ,\count_ones_reg[8]_i_1_n_5 ,\count_ones_reg[8]_i_1_n_6 ,\count_ones_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\count_ones_reg[8]_i_1_n_8 ,\count_ones_reg[8]_i_1_n_9 ,\count_ones_reg[8]_i_1_n_10 ,\count_ones_reg[8]_i_1_n_11 ,\count_ones_reg[8]_i_1_n_12 ,\count_ones_reg[8]_i_1_n_13 ,\count_ones_reg[8]_i_1_n_14 ,\count_ones_reg[8]_i_1_n_15 }),
        .S({\count_ones[8]_i_2_n_0 ,\count_ones[8]_i_3_n_0 ,\count_ones[8]_i_4_n_0 ,\count_ones[8]_i_5_n_0 ,\count_ones[8]_i_6_n_0 ,\count_ones[8]_i_7_n_0 ,\count_ones[8]_i_8_n_0 ,\count_ones[8]_i_9_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \count_ones_reg[9] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_ones_reg[8]_i_1_n_14 ),
        .Q(count_ones_reg[9]));
  LUT4 #(
    .INIT(16'h0004)) 
    \count_zeros[0]_i_10 
       (.I0(count_zeros_reg[0]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_2 
       (.I0(count_zeros_reg[0]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_3 
       (.I0(count_zeros_reg[7]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_4 
       (.I0(count_zeros_reg[6]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_5 
       (.I0(count_zeros_reg[5]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_6 
       (.I0(count_zeros_reg[4]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_7 
       (.I0(count_zeros_reg[3]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_8 
       (.I0(count_zeros_reg[2]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[0]_i_9 
       (.I0(count_zeros_reg[1]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[0]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[16]_i_2 
       (.I0(count_zeros_reg[16]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[16]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_2 
       (.I0(count_zeros_reg[15]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_3 
       (.I0(count_zeros_reg[14]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_4 
       (.I0(count_zeros_reg[13]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_5 
       (.I0(count_zeros_reg[12]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_6 
       (.I0(count_zeros_reg[11]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_7 
       (.I0(count_zeros_reg[10]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_8 
       (.I0(count_zeros_reg[9]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \count_zeros[8]_i_9 
       (.I0(count_zeros_reg[8]),
        .I1(ct_state[1]),
        .I2(ct_state[0]),
        .I3(ct_state[2]),
        .O(\count_zeros[8]_i_9_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[0] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_15 ),
        .Q(count_zeros_reg[0]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \count_zeros_reg[0]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\count_zeros_reg[0]_i_1_n_0 ,\count_zeros_reg[0]_i_1_n_1 ,\count_zeros_reg[0]_i_1_n_2 ,\count_zeros_reg[0]_i_1_n_3 ,\count_zeros_reg[0]_i_1_n_4 ,\count_zeros_reg[0]_i_1_n_5 ,\count_zeros_reg[0]_i_1_n_6 ,\count_zeros_reg[0]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\count_zeros[0]_i_2_n_0 }),
        .O({\count_zeros_reg[0]_i_1_n_8 ,\count_zeros_reg[0]_i_1_n_9 ,\count_zeros_reg[0]_i_1_n_10 ,\count_zeros_reg[0]_i_1_n_11 ,\count_zeros_reg[0]_i_1_n_12 ,\count_zeros_reg[0]_i_1_n_13 ,\count_zeros_reg[0]_i_1_n_14 ,\count_zeros_reg[0]_i_1_n_15 }),
        .S({\count_zeros[0]_i_3_n_0 ,\count_zeros[0]_i_4_n_0 ,\count_zeros[0]_i_5_n_0 ,\count_zeros[0]_i_6_n_0 ,\count_zeros[0]_i_7_n_0 ,\count_zeros[0]_i_8_n_0 ,\count_zeros[0]_i_9_n_0 ,\count_zeros[0]_i_10_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[10] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_13 ),
        .Q(count_zeros_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[11] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_12 ),
        .Q(count_zeros_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[12] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_11 ),
        .Q(count_zeros_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[13] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_10 ),
        .Q(count_zeros_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[14] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_9 ),
        .Q(count_zeros_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[15] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_8 ),
        .Q(count_zeros_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[16] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[16]_i_1_n_15 ),
        .Q(count_zeros_reg[16]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \count_zeros_reg[16]_i_1 
       (.CI(\count_zeros_reg[8]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO(\NLW_count_zeros_reg[16]_i_1_CO_UNCONNECTED [7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_count_zeros_reg[16]_i_1_O_UNCONNECTED [7:1],\count_zeros_reg[16]_i_1_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\count_zeros[16]_i_2_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[1] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_14 ),
        .Q(count_zeros_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[2] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_13 ),
        .Q(count_zeros_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[3] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_12 ),
        .Q(count_zeros_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[4] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_11 ),
        .Q(count_zeros_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[5] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_10 ),
        .Q(count_zeros_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[6] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_9 ),
        .Q(count_zeros_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[7] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[0]_i_1_n_8 ),
        .Q(count_zeros_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[8] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_15 ),
        .Q(count_zeros_reg[8]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \count_zeros_reg[8]_i_1 
       (.CI(\count_zeros_reg[0]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\count_zeros_reg[8]_i_1_n_0 ,\count_zeros_reg[8]_i_1_n_1 ,\count_zeros_reg[8]_i_1_n_2 ,\count_zeros_reg[8]_i_1_n_3 ,\count_zeros_reg[8]_i_1_n_4 ,\count_zeros_reg[8]_i_1_n_5 ,\count_zeros_reg[8]_i_1_n_6 ,\count_zeros_reg[8]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\count_zeros_reg[8]_i_1_n_8 ,\count_zeros_reg[8]_i_1_n_9 ,\count_zeros_reg[8]_i_1_n_10 ,\count_zeros_reg[8]_i_1_n_11 ,\count_zeros_reg[8]_i_1_n_12 ,\count_zeros_reg[8]_i_1_n_13 ,\count_zeros_reg[8]_i_1_n_14 ,\count_zeros_reg[8]_i_1_n_15 }),
        .S({\count_zeros[8]_i_2_n_0 ,\count_zeros[8]_i_3_n_0 ,\count_zeros[8]_i_4_n_0 ,\count_zeros[8]_i_5_n_0 ,\count_zeros[8]_i_6_n_0 ,\count_zeros[8]_i_7_n_0 ,\count_zeros[8]_i_8_n_0 ,\count_zeros[8]_i_9_n_0 }));
  FDCE #(
    .INIT(1'b0)) 
    \count_zeros_reg[9] 
       (.C(clk_i),
        .CE(count_ones),
        .CLR(rst_i),
        .D(\count_zeros_reg[8]_i_1_n_14 ),
        .Q(count_zeros_reg[9]));
  LUT6 #(
    .INIT(64'hFDDFFDD3FDDFFDDF)) 
    \ct_state[0]_i_1 
       (.I0(ce_i_d_reg_0),
        .I1(ct_state[0]),
        .I2(ct_state[2]),
        .I3(ct_state[1]),
        .I4(ce_i_d2),
        .I5(ce_i_d),
        .O(nxt_state[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF4400F444)) 
    \ct_state[1]_i_1 
       (.I0(load),
        .I1(ce_i_d_reg_0),
        .I2(\ct_state[2]_i_3_n_0 ),
        .I3(data_i_d2),
        .I4(data_i_d),
        .I5(\ct_state[1]_i_2_n_0 ),
        .O(nxt_state[1]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \ct_state[1]_i_2 
       (.I0(ce_i_d2),
        .I1(ce_i_d),
        .I2(ct_state[0]),
        .I3(out),
        .I4(ct_state[2]),
        .I5(ct_state[1]),
        .O(\ct_state[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F400F0)) 
    \ct_state[2]_i_1 
       (.I0(load),
        .I1(ce_i_d_reg_0),
        .I2(\ct_state[2]_i_3_n_0 ),
        .I3(data_i_d2),
        .I4(data_i_d),
        .I5(\ct_state[2]_i_4_n_0 ),
        .O(nxt_state[2]));
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \ct_state[2]_i_2 
       (.I0(ct_state[2]),
        .I1(ct_state[0]),
        .I2(ct_state[1]),
        .O(load));
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \ct_state[2]_i_3 
       (.I0(ct_state[0]),
        .I1(ce_i_d_reg_0),
        .I2(ct_state[1]),
        .I3(ct_state[2]),
        .O(\ct_state[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \ct_state[2]_i_4 
       (.I0(ce_i_d2),
        .I1(ce_i_d),
        .I2(ct_state[0]),
        .I3(out),
        .I4(ct_state[2]),
        .I5(ct_state[1]),
        .O(\ct_state[2]_i_4_n_0 ));
  (* FSM_ENCODED_STATES = "idle:001,cnt1:100,cnt0:010" *) 
  FDPE #(
    .INIT(1'b1)) 
    \ct_state_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(nxt_state[0]),
        .PRE(rst_i),
        .Q(ct_state[0]));
  (* FSM_ENCODED_STATES = "idle:001,cnt1:100,cnt0:010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \ct_state_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(nxt_state[1]),
        .Q(ct_state[1]));
  (* FSM_ENCODED_STATES = "idle:001,cnt1:100,cnt0:010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \ct_state_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(nxt_state[2]),
        .Q(ct_state[2]));
  FDCE #(
    .INIT(1'b0)) 
    data_i_d2_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(data_i_d),
        .Q(data_i_d2));
  FDCE #(
    .INIT(1'b0)) 
    data_i_d_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(out),
        .Q(data_i_d));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry__0_i_1
       (.I0(count_zeros_reg[16]),
        .O(i__carry__0_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry__0_i_1__0
       (.I0(count_ones_reg[16]),
        .O(i__carry__0_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry__0_i_1__1
       (.I0(count_zeros_reg[16]),
        .O(i__carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_1
       (.I0(count_zeros_reg[14]),
        .I1(count_zeros_reg[15]),
        .O(i__carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_10
       (.I0(count_ones_reg[6]),
        .I1(count_ones_reg[7]),
        .O(i__carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_10__0
       (.I0(count_zeros_reg[10]),
        .I1(count_zeros_reg[11]),
        .O(i__carry_i_10__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_10__1
       (.I0(count_zeros_reg[6]),
        .I1(count_zeros_reg[7]),
        .O(i__carry_i_10__1_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_10__4
       (.I0(count_zeros_reg[11]),
        .I1(count_zeros_reg[10]),
        .O(i__carry_i_10__4_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_11__0
       (.I0(count_zeros_reg[4]),
        .I1(count_zeros_reg[5]),
        .O(i__carry_i_11__0_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_11__1
       (.I0(count_zeros_reg[8]),
        .I1(count_zeros_reg[9]),
        .O(i__carry_i_11__1_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_11__2
       (.I0(count_zeros_reg[8]),
        .I1(count_zeros_reg[9]),
        .O(i__carry_i_11__2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_11__3
       (.I0(count_ones_reg[4]),
        .I1(count_ones_reg[5]),
        .O(i__carry_i_11__3_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_12
       (.I0(count_zeros_reg[6]),
        .I1(count_zeros_reg[7]),
        .O(i__carry_i_12_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_12__1
       (.I0(count_zeros_reg[7]),
        .I1(count_zeros_reg[6]),
        .O(i__carry_i_12__1_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_12__2
       (.I0(count_ones_reg[2]),
        .I1(count_ones_reg[3]),
        .O(i__carry_i_12__2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_12__3
       (.I0(count_zeros_reg[2]),
        .I1(count_zeros_reg[3]),
        .O(i__carry_i_12__3_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_13__0
       (.I0(count_zeros_reg[5]),
        .I1(count_zeros_reg[4]),
        .O(i__carry_i_13__0_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_13__1
       (.I0(count_zeros_reg[4]),
        .I1(count_zeros_reg[5]),
        .O(i__carry_i_13__1_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_13__2
       (.I0(count_ones_reg[0]),
        .I1(count_ones_reg[1]),
        .O(i__carry_i_13__2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_13__3
       (.I0(count_zeros_reg[0]),
        .I1(count_zeros_reg[1]),
        .O(i__carry_i_13__3_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_14__0
       (.I0(count_zeros_reg[3]),
        .I1(count_zeros_reg[2]),
        .O(i__carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_14__1
       (.I0(count_zeros_reg[2]),
        .I1(count_zeros_reg[3]),
        .O(i__carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_15__0
       (.I0(count_zeros_reg[0]),
        .I1(count_zeros_reg[1]),
        .O(i__carry_i_15__0_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_15__1
       (.I0(count_zeros_reg[0]),
        .I1(count_zeros_reg[1]),
        .O(i__carry_i_15__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_1__0
       (.I0(count_zeros_reg[14]),
        .I1(count_zeros_reg[15]),
        .O(i__carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_1__1
       (.I0(count_ones_reg[14]),
        .I1(count_ones_reg[15]),
        .O(i__carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    i__carry_i_1__4
       (.I0(count_zeros_reg[14]),
        .I1(count_zeros_reg[15]),
        .O(i__carry_i_1__4_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_2
       (.I0(count_ones_reg[12]),
        .I1(count_ones_reg[13]),
        .O(i__carry_i_2_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_2__0
       (.I0(count_zeros_reg[12]),
        .I1(count_zeros_reg[13]),
        .O(i__carry_i_2__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_2__1
       (.I0(count_zeros_reg[10]),
        .I1(count_zeros_reg[11]),
        .O(i__carry_i_2__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    i__carry_i_2__4
       (.I0(count_zeros_reg[12]),
        .I1(count_zeros_reg[13]),
        .O(i__carry_i_2__4_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_3
       (.I0(count_zeros_reg[8]),
        .I1(count_zeros_reg[9]),
        .O(i__carry_i_3_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_3__0
       (.I0(count_ones_reg[8]),
        .I1(count_ones_reg[9]),
        .O(i__carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_3__1
       (.I0(count_zeros_reg[8]),
        .I1(count_zeros_reg[9]),
        .O(i__carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    i__carry_i_3__4
       (.I0(count_zeros_reg[10]),
        .I1(count_zeros_reg[11]),
        .O(i__carry_i_3__4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_4
       (.I0(count_zeros_reg[6]),
        .I1(count_zeros_reg[7]),
        .O(i__carry_i_4_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_4__0
       (.I0(count_ones_reg[2]),
        .I1(count_ones_reg[3]),
        .O(i__carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_4__1
       (.I0(count_zeros_reg[2]),
        .I1(count_zeros_reg[3]),
        .O(i__carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_4__4
       (.I0(count_zeros_reg[8]),
        .I1(count_zeros_reg[9]),
        .O(i__carry_i_4__4_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_5
       (.I0(count_zeros_reg[4]),
        .I1(count_zeros_reg[5]),
        .O(i__carry_i_5_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_5__0
       (.I0(count_ones_reg[0]),
        .I1(count_ones_reg[1]),
        .O(i__carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_5__1
       (.I0(count_zeros_reg[0]),
        .I1(count_zeros_reg[1]),
        .O(i__carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    i__carry_i_5__4
       (.I0(count_zeros_reg[6]),
        .I1(count_zeros_reg[7]),
        .O(i__carry_i_5__4_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_6
       (.I0(count_zeros_reg[5]),
        .O(i__carry_i_6_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_6__0
       (.I0(count_zeros_reg[2]),
        .I1(count_zeros_reg[3]),
        .O(i__carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_6__3
       (.I0(count_ones_reg[15]),
        .I1(count_ones_reg[14]),
        .O(i__carry_i_6__3_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_6__4
       (.I0(count_zeros_reg[15]),
        .I1(count_zeros_reg[14]),
        .O(i__carry_i_6__4_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    i__carry_i_7
       (.I0(count_zeros_reg[3]),
        .O(i__carry_i_7_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    i__carry_i_7__0
       (.I0(count_zeros_reg[0]),
        .I1(count_zeros_reg[1]),
        .O(i__carry_i_7__0_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_7__3
       (.I0(count_ones_reg[12]),
        .I1(count_ones_reg[13]),
        .O(i__carry_i_7__3_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_7__4
       (.I0(count_zeros_reg[12]),
        .I1(count_zeros_reg[13]),
        .O(i__carry_i_7__4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_8
       (.I0(count_zeros_reg[14]),
        .I1(count_zeros_reg[15]),
        .O(i__carry_i_8_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_8__2
       (.I0(count_ones_reg[10]),
        .I1(count_ones_reg[11]),
        .O(i__carry_i_8__2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    i__carry_i_8__3
       (.I0(count_zeros_reg[10]),
        .I1(count_zeros_reg[11]),
        .O(i__carry_i_8__3_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_8__4
       (.I0(count_zeros_reg[14]),
        .I1(count_zeros_reg[15]),
        .O(i__carry_i_8__4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_9
       (.I0(count_zeros_reg[12]),
        .I1(count_zeros_reg[13]),
        .O(i__carry_i_9_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    i__carry_i_9__0
       (.I0(count_zeros_reg[12]),
        .I1(count_zeros_reg[13]),
        .O(i__carry_i_9__0_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_9__3
       (.I0(count_ones_reg[8]),
        .I1(count_ones_reg[9]),
        .O(i__carry_i_9__3_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    i__carry_i_9__4
       (.I0(count_zeros_reg[8]),
        .I1(count_zeros_reg[9]),
        .O(i__carry_i_9__4_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    q_o0_carry
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({q_o0_carry_n_0,q_o0_carry_n_1,q_o0_carry_n_2,q_o0_carry_n_3,q_o0_carry_n_4,q_o0_carry_n_5,q_o0_carry_n_6,q_o0_carry_n_7}),
        .DI({q_o0_carry_i_1_n_0,1'b0,q_o0_carry_i_2_n_0,q_o0_carry_i_3_n_0,q_o0_carry_i_4_n_0,q_o0_carry_i_5_n_0,q_o0_carry_i_6_n_0,q_o0_carry_i_7_n_0}),
        .O(NLW_q_o0_carry_O_UNCONNECTED[7:0]),
        .S({q_o0_carry_i_8_n_0,q_o0_carry_i_9_n_0,q_o0_carry_i_10_n_0,q_o0_carry_i_11_n_0,q_o0_carry_i_12_n_0,q_o0_carry_i_13_n_0,q_o0_carry_i_14_n_0,q_o0_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    q_o0_carry__0
       (.CI(q_o0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_q_o0_carry__0_CO_UNCONNECTED[7:1],double_one}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(NLW_q_o0_carry__0_O_UNCONNECTED[7:0]),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,count_ones_reg[16]}));
  LUT2 #(
    .INIT(4'hE)) 
    q_o0_carry_i_1
       (.I0(count_ones_reg[14]),
        .I1(count_ones_reg[15]),
        .O(q_o0_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    q_o0_carry_i_10
       (.I0(count_ones_reg[11]),
        .I1(count_ones_reg[10]),
        .O(q_o0_carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o0_carry_i_11
       (.I0(count_ones_reg[8]),
        .I1(count_ones_reg[9]),
        .O(q_o0_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    q_o0_carry_i_12
       (.I0(count_ones_reg[7]),
        .I1(count_ones_reg[6]),
        .O(q_o0_carry_i_12_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o0_carry_i_13
       (.I0(count_ones_reg[4]),
        .I1(count_ones_reg[5]),
        .O(q_o0_carry_i_13_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o0_carry_i_14
       (.I0(count_ones_reg[2]),
        .I1(count_ones_reg[3]),
        .O(q_o0_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o0_carry_i_15
       (.I0(count_ones_reg[0]),
        .I1(count_ones_reg[1]),
        .O(q_o0_carry_i_15_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o0_carry_i_2
       (.I0(count_ones_reg[10]),
        .I1(count_ones_reg[11]),
        .O(q_o0_carry_i_2_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    q_o0_carry_i_3
       (.I0(count_ones_reg[8]),
        .I1(count_ones_reg[9]),
        .O(q_o0_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o0_carry_i_4
       (.I0(count_ones_reg[6]),
        .I1(count_ones_reg[7]),
        .O(q_o0_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    q_o0_carry_i_5
       (.I0(count_ones_reg[4]),
        .I1(count_ones_reg[5]),
        .O(q_o0_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    q_o0_carry_i_6
       (.I0(count_ones_reg[2]),
        .I1(count_ones_reg[3]),
        .O(q_o0_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    q_o0_carry_i_7
       (.I0(count_ones_reg[0]),
        .I1(count_ones_reg[1]),
        .O(q_o0_carry_i_7_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o0_carry_i_8
       (.I0(count_ones_reg[14]),
        .I1(count_ones_reg[15]),
        .O(q_o0_carry_i_8_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o0_carry_i_9
       (.I0(count_ones_reg[12]),
        .I1(count_ones_reg[13]),
        .O(q_o0_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o0_inferred__0/i__carry 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\q_o0_inferred__0/i__carry_n_0 ,\q_o0_inferred__0/i__carry_n_1 ,\q_o0_inferred__0/i__carry_n_2 ,\q_o0_inferred__0/i__carry_n_3 ,\q_o0_inferred__0/i__carry_n_4 ,\q_o0_inferred__0/i__carry_n_5 ,\q_o0_inferred__0/i__carry_n_6 ,\q_o0_inferred__0/i__carry_n_7 }),
        .DI({i__carry_i_1_n_0,1'b0,i__carry_i_2__1_n_0,i__carry_i_3_n_0,i__carry_i_4_n_0,i__carry_i_5_n_0,i__carry_i_6__0_n_0,i__carry_i_7__0_n_0}),
        .O(\NLW_q_o0_inferred__0/i__carry_O_UNCONNECTED [7:0]),
        .S({i__carry_i_8__4_n_0,i__carry_i_9_n_0,i__carry_i_10__4_n_0,i__carry_i_11__2_n_0,i__carry_i_12__1_n_0,i__carry_i_13__1_n_0,i__carry_i_14__1_n_0,i__carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o0_inferred__0/i__carry__0 
       (.CI(\q_o0_inferred__0/i__carry_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_q_o0_inferred__0/i__carry__0_CO_UNCONNECTED [7:1],\count_zeros_reg[16]_1 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(\NLW_q_o0_inferred__0/i__carry__0_O_UNCONNECTED [7:0]),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,count_zeros_reg[16]}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    q_o1_carry
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({q_o1_carry_n_0,q_o1_carry_n_1,q_o1_carry_n_2,q_o1_carry_n_3,q_o1_carry_n_4,q_o1_carry_n_5,q_o1_carry_n_6,q_o1_carry_n_7}),
        .DI({q_o1_carry_i_1_n_0,q_o1_carry_i_2_n_0,q_o1_carry_i_3_n_0,q_o1_carry_i_4_n_0,q_o1_carry_i_5_n_0,q_o1_carry_i_6_n_0,q_o1_carry_i_7_n_0,1'b0}),
        .O(NLW_q_o1_carry_O_UNCONNECTED[7:0]),
        .S({q_o1_carry_i_8_n_0,q_o1_carry_i_9_n_0,q_o1_carry_i_10_n_0,q_o1_carry_i_11_n_0,q_o1_carry_i_12_n_0,q_o1_carry_i_13_n_0,q_o1_carry_i_14_n_0,q_o1_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    q_o1_carry__0
       (.CI(q_o1_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_q_o1_carry__0_CO_UNCONNECTED[7:1],q_o1}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(NLW_q_o1_carry__0_O_UNCONNECTED[7:0]),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,q_o1_carry__0_i_1_n_0}));
  LUT1 #(
    .INIT(2'h1)) 
    q_o1_carry__0_i_1
       (.I0(count_ones_reg[16]),
        .O(q_o1_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    q_o1_carry_i_1
       (.I0(count_ones_reg[14]),
        .I1(count_ones_reg[15]),
        .O(q_o1_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o1_carry_i_10
       (.I0(count_ones_reg[10]),
        .I1(count_ones_reg[11]),
        .O(q_o1_carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    q_o1_carry_i_11
       (.I0(count_ones_reg[8]),
        .I1(count_ones_reg[9]),
        .O(q_o1_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o1_carry_i_12
       (.I0(count_ones_reg[6]),
        .I1(count_ones_reg[7]),
        .O(q_o1_carry_i_12_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    q_o1_carry_i_13
       (.I0(count_ones_reg[5]),
        .I1(count_ones_reg[4]),
        .O(q_o1_carry_i_13_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    q_o1_carry_i_14
       (.I0(count_ones_reg[3]),
        .I1(count_ones_reg[2]),
        .O(q_o1_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o1_carry_i_15
       (.I0(count_ones_reg[0]),
        .I1(count_ones_reg[1]),
        .O(q_o1_carry_i_15_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    q_o1_carry_i_2
       (.I0(count_ones_reg[12]),
        .I1(count_ones_reg[13]),
        .O(q_o1_carry_i_2_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    q_o1_carry_i_3
       (.I0(count_ones_reg[10]),
        .I1(count_ones_reg[11]),
        .O(q_o1_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    q_o1_carry_i_4
       (.I0(count_ones_reg[8]),
        .I1(count_ones_reg[9]),
        .O(q_o1_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    q_o1_carry_i_5
       (.I0(count_ones_reg[6]),
        .I1(count_ones_reg[7]),
        .O(q_o1_carry_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    q_o1_carry_i_6
       (.I0(count_ones_reg[5]),
        .O(q_o1_carry_i_6_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    q_o1_carry_i_7
       (.I0(count_ones_reg[3]),
        .O(q_o1_carry_i_7_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o1_carry_i_8
       (.I0(count_ones_reg[14]),
        .I1(count_ones_reg[15]),
        .O(q_o1_carry_i_8_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    q_o1_carry_i_9
       (.I0(count_ones_reg[12]),
        .I1(count_ones_reg[13]),
        .O(q_o1_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o1_inferred__0/i__carry 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\q_o1_inferred__0/i__carry_n_0 ,\q_o1_inferred__0/i__carry_n_1 ,\q_o1_inferred__0/i__carry_n_2 ,\q_o1_inferred__0/i__carry_n_3 ,\q_o1_inferred__0/i__carry_n_4 ,\q_o1_inferred__0/i__carry_n_5 ,\q_o1_inferred__0/i__carry_n_6 ,\q_o1_inferred__0/i__carry_n_7 }),
        .DI({i__carry_i_1__1_n_0,i__carry_i_2_n_0,count_ones_reg[11],i__carry_i_3__0_n_0,1'b0,count_ones_reg[5],i__carry_i_4__0_n_0,i__carry_i_5__0_n_0}),
        .O(\NLW_q_o1_inferred__0/i__carry_O_UNCONNECTED [7:0]),
        .S({i__carry_i_6__3_n_0,i__carry_i_7__3_n_0,i__carry_i_8__2_n_0,i__carry_i_9__3_n_0,i__carry_i_10_n_0,i__carry_i_11__3_n_0,i__carry_i_12__2_n_0,i__carry_i_13__2_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o1_inferred__0/i__carry__0 
       (.CI(\q_o1_inferred__0/i__carry_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_q_o1_inferred__0/i__carry__0_CO_UNCONNECTED [7:1],q_o10_in}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,count_ones_reg[16]}),
        .O(\NLW_q_o1_inferred__0/i__carry__0_O_UNCONNECTED [7:0]),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,i__carry__0_i_1__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o1_inferred__1/i__carry 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\q_o1_inferred__1/i__carry_n_0 ,\q_o1_inferred__1/i__carry_n_1 ,\q_o1_inferred__1/i__carry_n_2 ,\q_o1_inferred__1/i__carry_n_3 ,\q_o1_inferred__1/i__carry_n_4 ,\q_o1_inferred__1/i__carry_n_5 ,\q_o1_inferred__1/i__carry_n_6 ,\q_o1_inferred__1/i__carry_n_7 }),
        .DI({i__carry_i_1__4_n_0,i__carry_i_2__4_n_0,i__carry_i_3__4_n_0,i__carry_i_4__4_n_0,i__carry_i_5__4_n_0,i__carry_i_6_n_0,i__carry_i_7_n_0,1'b0}),
        .O(\NLW_q_o1_inferred__1/i__carry_O_UNCONNECTED [7:0]),
        .S({i__carry_i_8_n_0,i__carry_i_9__0_n_0,i__carry_i_10__0_n_0,i__carry_i_11__1_n_0,i__carry_i_12_n_0,i__carry_i_13__0_n_0,i__carry_i_14__0_n_0,i__carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o1_inferred__1/i__carry__0 
       (.CI(\q_o1_inferred__1/i__carry_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_q_o1_inferred__1/i__carry__0_CO_UNCONNECTED [7:1],CO}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(\NLW_q_o1_inferred__1/i__carry__0_O_UNCONNECTED [7:0]),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,i__carry__0_i_1__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o1_inferred__2/i__carry 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\q_o1_inferred__2/i__carry_n_0 ,\q_o1_inferred__2/i__carry_n_1 ,\q_o1_inferred__2/i__carry_n_2 ,\q_o1_inferred__2/i__carry_n_3 ,\q_o1_inferred__2/i__carry_n_4 ,\q_o1_inferred__2/i__carry_n_5 ,\q_o1_inferred__2/i__carry_n_6 ,\q_o1_inferred__2/i__carry_n_7 }),
        .DI({i__carry_i_1__0_n_0,i__carry_i_2__0_n_0,count_zeros_reg[11],i__carry_i_3__1_n_0,1'b0,count_zeros_reg[5],i__carry_i_4__1_n_0,i__carry_i_5__1_n_0}),
        .O(\NLW_q_o1_inferred__2/i__carry_O_UNCONNECTED [7:0]),
        .S({i__carry_i_6__4_n_0,i__carry_i_7__4_n_0,i__carry_i_8__3_n_0,i__carry_i_9__4_n_0,i__carry_i_10__1_n_0,i__carry_i_11__0_n_0,i__carry_i_12__3_n_0,i__carry_i_13__3_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \q_o1_inferred__2/i__carry__0 
       (.CI(\q_o1_inferred__2/i__carry_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_q_o1_inferred__2/i__carry__0_CO_UNCONNECTED [7:1],\count_zeros_reg[16]_0 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,count_zeros_reg[16]}),
        .O(\NLW_q_o1_inferred__2/i__carry__0_O_UNCONNECTED [7:0]),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,i__carry__0_i_1_n_0}));
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT2 #(
    .INIT(4'h2)) 
    recieved_debug_inferred_i_1
       (.I0(\count_zeros_reg[16]_1 ),
        .I1(rst_i),
        .O(in0[3]));
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'h08)) 
    recieved_debug_inferred_i_2
       (.I0(CO),
        .I1(\count_zeros_reg[16]_0 ),
        .I2(rst_i),
        .O(in0[2]));
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT2 #(
    .INIT(4'h2)) 
    recieved_debug_inferred_i_3
       (.I0(double_one),
        .I1(rst_i),
        .O(in0[1]));
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'h08)) 
    recieved_debug_inferred_i_4
       (.I0(q_o1),
        .I1(q_o10_in),
        .I2(rst_i),
        .O(in0[0]));
endmodule

(* ORIG_REF_NAME = "waitForStart" *) 
module switch_elements_waitForStart
   (waitforstart_rdy,
    clk_i,
    rst_i,
    out);
  output waitforstart_rdy;
  input clk_i;
  input rst_i;
  input out;

  wire clk_i;
  wire [31:0]counter;
  wire counter0_carry__0_n_0;
  wire counter0_carry__0_n_1;
  wire counter0_carry__0_n_10;
  wire counter0_carry__0_n_11;
  wire counter0_carry__0_n_12;
  wire counter0_carry__0_n_13;
  wire counter0_carry__0_n_14;
  wire counter0_carry__0_n_15;
  wire counter0_carry__0_n_2;
  wire counter0_carry__0_n_3;
  wire counter0_carry__0_n_4;
  wire counter0_carry__0_n_5;
  wire counter0_carry__0_n_6;
  wire counter0_carry__0_n_7;
  wire counter0_carry__0_n_8;
  wire counter0_carry__0_n_9;
  wire counter0_carry__1_n_0;
  wire counter0_carry__1_n_1;
  wire counter0_carry__1_n_10;
  wire counter0_carry__1_n_11;
  wire counter0_carry__1_n_12;
  wire counter0_carry__1_n_13;
  wire counter0_carry__1_n_14;
  wire counter0_carry__1_n_15;
  wire counter0_carry__1_n_2;
  wire counter0_carry__1_n_3;
  wire counter0_carry__1_n_4;
  wire counter0_carry__1_n_5;
  wire counter0_carry__1_n_6;
  wire counter0_carry__1_n_7;
  wire counter0_carry__1_n_8;
  wire counter0_carry__1_n_9;
  wire counter0_carry__2_n_10;
  wire counter0_carry__2_n_11;
  wire counter0_carry__2_n_12;
  wire counter0_carry__2_n_13;
  wire counter0_carry__2_n_14;
  wire counter0_carry__2_n_15;
  wire counter0_carry__2_n_2;
  wire counter0_carry__2_n_3;
  wire counter0_carry__2_n_4;
  wire counter0_carry__2_n_5;
  wire counter0_carry__2_n_6;
  wire counter0_carry__2_n_7;
  wire counter0_carry__2_n_9;
  wire counter0_carry_n_0;
  wire counter0_carry_n_1;
  wire counter0_carry_n_10;
  wire counter0_carry_n_11;
  wire counter0_carry_n_12;
  wire counter0_carry_n_13;
  wire counter0_carry_n_14;
  wire counter0_carry_n_15;
  wire counter0_carry_n_2;
  wire counter0_carry_n_3;
  wire counter0_carry_n_4;
  wire counter0_carry_n_5;
  wire counter0_carry_n_6;
  wire counter0_carry_n_7;
  wire counter0_carry_n_8;
  wire counter0_carry_n_9;
  wire \counter_reg_n_0_[0] ;
  wire \counter_reg_n_0_[10] ;
  wire \counter_reg_n_0_[11] ;
  wire \counter_reg_n_0_[12] ;
  wire \counter_reg_n_0_[13] ;
  wire \counter_reg_n_0_[14] ;
  wire \counter_reg_n_0_[15] ;
  wire \counter_reg_n_0_[16] ;
  wire \counter_reg_n_0_[17] ;
  wire \counter_reg_n_0_[18] ;
  wire \counter_reg_n_0_[19] ;
  wire \counter_reg_n_0_[1] ;
  wire \counter_reg_n_0_[20] ;
  wire \counter_reg_n_0_[21] ;
  wire \counter_reg_n_0_[22] ;
  wire \counter_reg_n_0_[23] ;
  wire \counter_reg_n_0_[24] ;
  wire \counter_reg_n_0_[25] ;
  wire \counter_reg_n_0_[26] ;
  wire \counter_reg_n_0_[27] ;
  wire \counter_reg_n_0_[28] ;
  wire \counter_reg_n_0_[29] ;
  wire \counter_reg_n_0_[2] ;
  wire \counter_reg_n_0_[30] ;
  wire \counter_reg_n_0_[31] ;
  wire \counter_reg_n_0_[3] ;
  wire \counter_reg_n_0_[4] ;
  wire \counter_reg_n_0_[5] ;
  wire \counter_reg_n_0_[6] ;
  wire \counter_reg_n_0_[7] ;
  wire \counter_reg_n_0_[8] ;
  wire \counter_reg_n_0_[9] ;
  wire lock;
  wire out;
  wire ready_o1_carry__0_i_10_n_0;
  wire ready_o1_carry__0_i_11_n_0;
  wire ready_o1_carry__0_i_12_n_0;
  wire ready_o1_carry__0_i_13_n_0;
  wire ready_o1_carry__0_i_14_n_0;
  wire ready_o1_carry__0_i_1_n_0;
  wire ready_o1_carry__0_i_2_n_0;
  wire ready_o1_carry__0_i_3_n_0;
  wire ready_o1_carry__0_i_4_n_0;
  wire ready_o1_carry__0_i_5_n_0;
  wire ready_o1_carry__0_i_6_n_0;
  wire ready_o1_carry__0_i_7_n_0;
  wire ready_o1_carry__0_i_8_n_0;
  wire ready_o1_carry__0_i_9_n_0;
  wire ready_o1_carry__0_n_1;
  wire ready_o1_carry__0_n_2;
  wire ready_o1_carry__0_n_3;
  wire ready_o1_carry__0_n_4;
  wire ready_o1_carry__0_n_5;
  wire ready_o1_carry__0_n_6;
  wire ready_o1_carry__0_n_7;
  wire ready_o1_carry_i_10_n_0;
  wire ready_o1_carry_i_11_n_0;
  wire ready_o1_carry_i_12_n_0;
  wire ready_o1_carry_i_13_n_0;
  wire ready_o1_carry_i_14_n_0;
  wire ready_o1_carry_i_15_n_0;
  wire ready_o1_carry_i_1_n_0;
  wire ready_o1_carry_i_2_n_0;
  wire ready_o1_carry_i_3_n_0;
  wire ready_o1_carry_i_4_n_0;
  wire ready_o1_carry_i_5_n_0;
  wire ready_o1_carry_i_6_n_0;
  wire ready_o1_carry_i_7_n_0;
  wire ready_o1_carry_i_8_n_0;
  wire ready_o1_carry_i_9_n_0;
  wire ready_o1_carry_n_0;
  wire ready_o1_carry_n_1;
  wire ready_o1_carry_n_2;
  wire ready_o1_carry_n_3;
  wire ready_o1_carry_n_4;
  wire ready_o1_carry_n_5;
  wire ready_o1_carry_n_6;
  wire ready_o1_carry_n_7;
  wire ready_o_i_1_n_0;
  wire rst_i;
  wire waitforstart_rdy;
  wire [7:6]NLW_counter0_carry__2_CO_UNCONNECTED;
  wire [7:7]NLW_counter0_carry__2_O_UNCONNECTED;
  wire [7:0]NLW_ready_o1_carry_O_UNCONNECTED;
  wire [7:7]NLW_ready_o1_carry__0_CO_UNCONNECTED;
  wire [7:0]NLW_ready_o1_carry__0_O_UNCONNECTED;

  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    counter0_carry
       (.CI(\counter_reg_n_0_[0] ),
        .CI_TOP(1'b0),
        .CO({counter0_carry_n_0,counter0_carry_n_1,counter0_carry_n_2,counter0_carry_n_3,counter0_carry_n_4,counter0_carry_n_5,counter0_carry_n_6,counter0_carry_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({counter0_carry_n_8,counter0_carry_n_9,counter0_carry_n_10,counter0_carry_n_11,counter0_carry_n_12,counter0_carry_n_13,counter0_carry_n_14,counter0_carry_n_15}),
        .S({\counter_reg_n_0_[8] ,\counter_reg_n_0_[7] ,\counter_reg_n_0_[6] ,\counter_reg_n_0_[5] ,\counter_reg_n_0_[4] ,\counter_reg_n_0_[3] ,\counter_reg_n_0_[2] ,\counter_reg_n_0_[1] }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    counter0_carry__0
       (.CI(counter0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({counter0_carry__0_n_0,counter0_carry__0_n_1,counter0_carry__0_n_2,counter0_carry__0_n_3,counter0_carry__0_n_4,counter0_carry__0_n_5,counter0_carry__0_n_6,counter0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({counter0_carry__0_n_8,counter0_carry__0_n_9,counter0_carry__0_n_10,counter0_carry__0_n_11,counter0_carry__0_n_12,counter0_carry__0_n_13,counter0_carry__0_n_14,counter0_carry__0_n_15}),
        .S({\counter_reg_n_0_[16] ,\counter_reg_n_0_[15] ,\counter_reg_n_0_[14] ,\counter_reg_n_0_[13] ,\counter_reg_n_0_[12] ,\counter_reg_n_0_[11] ,\counter_reg_n_0_[10] ,\counter_reg_n_0_[9] }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    counter0_carry__1
       (.CI(counter0_carry__0_n_0),
        .CI_TOP(1'b0),
        .CO({counter0_carry__1_n_0,counter0_carry__1_n_1,counter0_carry__1_n_2,counter0_carry__1_n_3,counter0_carry__1_n_4,counter0_carry__1_n_5,counter0_carry__1_n_6,counter0_carry__1_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({counter0_carry__1_n_8,counter0_carry__1_n_9,counter0_carry__1_n_10,counter0_carry__1_n_11,counter0_carry__1_n_12,counter0_carry__1_n_13,counter0_carry__1_n_14,counter0_carry__1_n_15}),
        .S({\counter_reg_n_0_[24] ,\counter_reg_n_0_[23] ,\counter_reg_n_0_[22] ,\counter_reg_n_0_[21] ,\counter_reg_n_0_[20] ,\counter_reg_n_0_[19] ,\counter_reg_n_0_[18] ,\counter_reg_n_0_[17] }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    counter0_carry__2
       (.CI(counter0_carry__1_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_counter0_carry__2_CO_UNCONNECTED[7:6],counter0_carry__2_n_2,counter0_carry__2_n_3,counter0_carry__2_n_4,counter0_carry__2_n_5,counter0_carry__2_n_6,counter0_carry__2_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_counter0_carry__2_O_UNCONNECTED[7],counter0_carry__2_n_9,counter0_carry__2_n_10,counter0_carry__2_n_11,counter0_carry__2_n_12,counter0_carry__2_n_13,counter0_carry__2_n_14,counter0_carry__2_n_15}),
        .S({1'b0,\counter_reg_n_0_[31] ,\counter_reg_n_0_[30] ,\counter_reg_n_0_[29] ,\counter_reg_n_0_[28] ,\counter_reg_n_0_[27] ,\counter_reg_n_0_[26] ,\counter_reg_n_0_[25] }));
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \counter[0]_i_1 
       (.I0(out),
        .I1(\counter_reg_n_0_[0] ),
        .O(counter[0]));
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[10]_i_1 
       (.I0(counter0_carry__0_n_14),
        .I1(out),
        .O(counter[10]));
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[11]_i_1 
       (.I0(counter0_carry__0_n_13),
        .I1(out),
        .O(counter[11]));
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[12]_i_1 
       (.I0(counter0_carry__0_n_12),
        .I1(out),
        .O(counter[12]));
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[13]_i_1 
       (.I0(counter0_carry__0_n_11),
        .I1(out),
        .O(counter[13]));
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[14]_i_1 
       (.I0(counter0_carry__0_n_10),
        .I1(out),
        .O(counter[14]));
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[15]_i_1 
       (.I0(counter0_carry__0_n_9),
        .I1(out),
        .O(counter[15]));
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[16]_i_1 
       (.I0(counter0_carry__0_n_8),
        .I1(out),
        .O(counter[16]));
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[17]_i_1 
       (.I0(counter0_carry__1_n_15),
        .I1(out),
        .O(counter[17]));
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[18]_i_1 
       (.I0(counter0_carry__1_n_14),
        .I1(out),
        .O(counter[18]));
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[19]_i_1 
       (.I0(counter0_carry__1_n_13),
        .I1(out),
        .O(counter[19]));
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[1]_i_1 
       (.I0(counter0_carry_n_15),
        .I1(out),
        .O(counter[1]));
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[20]_i_1 
       (.I0(counter0_carry__1_n_12),
        .I1(out),
        .O(counter[20]));
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[21]_i_1 
       (.I0(counter0_carry__1_n_11),
        .I1(out),
        .O(counter[21]));
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[22]_i_1 
       (.I0(counter0_carry__1_n_10),
        .I1(out),
        .O(counter[22]));
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[23]_i_1 
       (.I0(counter0_carry__1_n_9),
        .I1(out),
        .O(counter[23]));
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[24]_i_1 
       (.I0(counter0_carry__1_n_8),
        .I1(out),
        .O(counter[24]));
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[25]_i_1 
       (.I0(counter0_carry__2_n_15),
        .I1(out),
        .O(counter[25]));
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[26]_i_1 
       (.I0(counter0_carry__2_n_14),
        .I1(out),
        .O(counter[26]));
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[27]_i_1 
       (.I0(counter0_carry__2_n_13),
        .I1(out),
        .O(counter[27]));
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[28]_i_1 
       (.I0(counter0_carry__2_n_12),
        .I1(out),
        .O(counter[28]));
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[29]_i_1 
       (.I0(counter0_carry__2_n_11),
        .I1(out),
        .O(counter[29]));
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[2]_i_1 
       (.I0(counter0_carry_n_14),
        .I1(out),
        .O(counter[2]));
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[30]_i_1 
       (.I0(counter0_carry__2_n_10),
        .I1(out),
        .O(counter[30]));
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[31]_i_1 
       (.I0(counter0_carry__2_n_9),
        .I1(out),
        .O(counter[31]));
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[3]_i_1 
       (.I0(counter0_carry_n_13),
        .I1(out),
        .O(counter[3]));
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[4]_i_1 
       (.I0(counter0_carry_n_12),
        .I1(out),
        .O(counter[4]));
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[5]_i_1 
       (.I0(counter0_carry_n_11),
        .I1(out),
        .O(counter[5]));
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[6]_i_1 
       (.I0(counter0_carry_n_10),
        .I1(out),
        .O(counter[6]));
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[7]_i_1 
       (.I0(counter0_carry_n_9),
        .I1(out),
        .O(counter[7]));
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[8]_i_1 
       (.I0(counter0_carry_n_8),
        .I1(out),
        .O(counter[8]));
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \counter[9]_i_1 
       (.I0(counter0_carry__0_n_15),
        .I1(out),
        .O(counter[9]));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[0]),
        .Q(\counter_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[10]),
        .Q(\counter_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[11]),
        .Q(\counter_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[12]),
        .Q(\counter_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[13]),
        .Q(\counter_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[14]),
        .Q(\counter_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[15]),
        .Q(\counter_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[16]),
        .Q(\counter_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[17]),
        .Q(\counter_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[18]),
        .Q(\counter_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[19]),
        .Q(\counter_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[1]),
        .Q(\counter_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[20]),
        .Q(\counter_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[21]),
        .Q(\counter_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[22]),
        .Q(\counter_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[23]),
        .Q(\counter_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[24]),
        .Q(\counter_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[25]),
        .Q(\counter_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[26]),
        .Q(\counter_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[27]),
        .Q(\counter_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[28]),
        .Q(\counter_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[29]),
        .Q(\counter_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[2]),
        .Q(\counter_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[30]),
        .Q(\counter_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[31]),
        .Q(\counter_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[3]),
        .Q(\counter_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[4]),
        .Q(\counter_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[5]),
        .Q(\counter_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[6]),
        .Q(\counter_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[7]),
        .Q(\counter_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[8]),
        .Q(\counter_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \counter_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(counter[9]),
        .Q(\counter_reg_n_0_[9] ));
  FDCE #(
    .INIT(1'b0)) 
    lock_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(ready_o_i_1_n_0),
        .Q(lock));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    ready_o1_carry
       (.CI(ready_o1_carry_i_1_n_0),
        .CI_TOP(1'b0),
        .CO({ready_o1_carry_n_0,ready_o1_carry_n_1,ready_o1_carry_n_2,ready_o1_carry_n_3,ready_o1_carry_n_4,ready_o1_carry_n_5,ready_o1_carry_n_6,ready_o1_carry_n_7}),
        .DI({ready_o1_carry_i_2_n_0,1'b0,ready_o1_carry_i_3_n_0,ready_o1_carry_i_4_n_0,1'b0,ready_o1_carry_i_5_n_0,ready_o1_carry_i_6_n_0,ready_o1_carry_i_7_n_0}),
        .O(NLW_ready_o1_carry_O_UNCONNECTED[7:0]),
        .S({ready_o1_carry_i_8_n_0,ready_o1_carry_i_9_n_0,ready_o1_carry_i_10_n_0,ready_o1_carry_i_11_n_0,ready_o1_carry_i_12_n_0,ready_o1_carry_i_13_n_0,ready_o1_carry_i_14_n_0,ready_o1_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    ready_o1_carry__0
       (.CI(ready_o1_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_ready_o1_carry__0_CO_UNCONNECTED[7],ready_o1_carry__0_n_1,ready_o1_carry__0_n_2,ready_o1_carry__0_n_3,ready_o1_carry__0_n_4,ready_o1_carry__0_n_5,ready_o1_carry__0_n_6,ready_o1_carry__0_n_7}),
        .DI({1'b0,ready_o1_carry__0_i_1_n_0,ready_o1_carry__0_i_2_n_0,ready_o1_carry__0_i_3_n_0,ready_o1_carry__0_i_4_n_0,ready_o1_carry__0_i_5_n_0,ready_o1_carry__0_i_6_n_0,ready_o1_carry__0_i_7_n_0}),
        .O(NLW_ready_o1_carry__0_O_UNCONNECTED[7:0]),
        .S({1'b0,ready_o1_carry__0_i_8_n_0,ready_o1_carry__0_i_9_n_0,ready_o1_carry__0_i_10_n_0,ready_o1_carry__0_i_11_n_0,ready_o1_carry__0_i_12_n_0,ready_o1_carry__0_i_13_n_0,ready_o1_carry__0_i_14_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    ready_o1_carry__0_i_1
       (.I0(counter0_carry__2_n_9),
        .I1(out),
        .I2(counter0_carry__2_n_10),
        .O(ready_o1_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry__0_i_10
       (.I0(counter0_carry__2_n_13),
        .I1(counter0_carry__2_n_14),
        .I2(out),
        .O(ready_o1_carry__0_i_10_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry__0_i_11
       (.I0(counter0_carry__2_n_15),
        .I1(counter0_carry__1_n_8),
        .I2(out),
        .O(ready_o1_carry__0_i_11_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry__0_i_12
       (.I0(counter0_carry__1_n_9),
        .I1(counter0_carry__1_n_10),
        .I2(out),
        .O(ready_o1_carry__0_i_12_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry__0_i_13
       (.I0(counter0_carry__1_n_11),
        .I1(counter0_carry__1_n_12),
        .I2(out),
        .O(ready_o1_carry__0_i_13_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    ready_o1_carry__0_i_14
       (.I0(out),
        .I1(counter0_carry__1_n_13),
        .I2(counter0_carry__1_n_14),
        .O(ready_o1_carry__0_i_14_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry__0_i_2
       (.I0(out),
        .I1(counter0_carry__2_n_12),
        .I2(counter0_carry__2_n_11),
        .O(ready_o1_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry__0_i_3
       (.I0(out),
        .I1(counter0_carry__2_n_14),
        .I2(counter0_carry__2_n_13),
        .O(ready_o1_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry__0_i_4
       (.I0(out),
        .I1(counter0_carry__1_n_8),
        .I2(counter0_carry__2_n_15),
        .O(ready_o1_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry__0_i_5
       (.I0(out),
        .I1(counter0_carry__1_n_10),
        .I2(counter0_carry__1_n_9),
        .O(ready_o1_carry__0_i_5_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry__0_i_6
       (.I0(out),
        .I1(counter0_carry__1_n_12),
        .I2(counter0_carry__1_n_11),
        .O(ready_o1_carry__0_i_6_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ready_o1_carry__0_i_7
       (.I0(out),
        .I1(counter0_carry__1_n_13),
        .I2(counter0_carry__1_n_14),
        .O(ready_o1_carry__0_i_7_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry__0_i_8
       (.I0(counter0_carry__2_n_9),
        .I1(counter0_carry__2_n_10),
        .I2(out),
        .O(ready_o1_carry__0_i_8_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry__0_i_9
       (.I0(counter0_carry__2_n_11),
        .I1(counter0_carry__2_n_12),
        .I2(out),
        .O(ready_o1_carry__0_i_9_n_0));
  LUT3 #(
    .INIT(8'hD0)) 
    ready_o1_carry_i_1
       (.I0(\counter_reg_n_0_[0] ),
        .I1(counter0_carry_n_15),
        .I2(out),
        .O(ready_o1_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    ready_o1_carry_i_10
       (.I0(out),
        .I1(counter0_carry__0_n_11),
        .I2(counter0_carry__0_n_12),
        .O(ready_o1_carry_i_10_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    ready_o1_carry_i_11
       (.I0(out),
        .I1(counter0_carry__0_n_13),
        .I2(counter0_carry__0_n_14),
        .O(ready_o1_carry_i_11_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ready_o1_carry_i_12
       (.I0(out),
        .I1(counter0_carry__0_n_15),
        .I2(counter0_carry_n_8),
        .O(ready_o1_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry_i_13
       (.I0(counter0_carry_n_9),
        .I1(counter0_carry_n_10),
        .I2(out),
        .O(ready_o1_carry_i_13_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    ready_o1_carry_i_14
       (.I0(counter0_carry_n_11),
        .I1(out),
        .I2(counter0_carry_n_12),
        .O(ready_o1_carry_i_14_n_0));
  LUT3 #(
    .INIT(8'h1F)) 
    ready_o1_carry_i_15
       (.I0(counter0_carry_n_13),
        .I1(counter0_carry_n_14),
        .I2(out),
        .O(ready_o1_carry_i_15_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ready_o1_carry_i_2
       (.I0(counter0_carry__1_n_15),
        .I1(out),
        .O(ready_o1_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ready_o1_carry_i_3
       (.I0(out),
        .I1(counter0_carry__0_n_11),
        .I2(counter0_carry__0_n_12),
        .O(ready_o1_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ready_o1_carry_i_4
       (.I0(out),
        .I1(counter0_carry__0_n_13),
        .I2(counter0_carry__0_n_14),
        .O(ready_o1_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry_i_5
       (.I0(out),
        .I1(counter0_carry_n_10),
        .I2(counter0_carry_n_9),
        .O(ready_o1_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ready_o1_carry_i_6
       (.I0(counter0_carry_n_11),
        .I1(out),
        .O(ready_o1_carry_i_6_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    ready_o1_carry_i_7
       (.I0(out),
        .I1(counter0_carry_n_14),
        .I2(counter0_carry_n_13),
        .O(ready_o1_carry_i_7_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    ready_o1_carry_i_8
       (.I0(counter0_carry__1_n_15),
        .I1(out),
        .I2(counter0_carry__0_n_8),
        .O(ready_o1_carry_i_8_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ready_o1_carry_i_9
       (.I0(out),
        .I1(counter0_carry__0_n_9),
        .I2(counter0_carry__0_n_10),
        .O(ready_o1_carry_i_9_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ready_o_i_1
       (.I0(ready_o1_carry__0_n_1),
        .I1(lock),
        .O(ready_o_i_1_n_0));
  FDCE #(
    .INIT(1'b0)) 
    ready_o_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(ready_o_i_1_n_0),
        .Q(waitforstart_rdy));
endmodule
`ifndef GLBL
`define GLBL
`timescale  1 ps / 1 ps

module glbl ();

    parameter ROC_WIDTH = 100000;
    parameter TOC_WIDTH = 0;

//--------   STARTUP Globals --------------
    wire GSR;
    wire GTS;
    wire GWE;
    wire PRLD;
    tri1 p_up_tmp;
    tri (weak1, strong0) PLL_LOCKG = p_up_tmp;

    wire PROGB_GLBL;
    wire CCLKO_GLBL;
    wire FCSBO_GLBL;
    wire [3:0] DO_GLBL;
    wire [3:0] DI_GLBL;
   
    reg GSR_int;
    reg GTS_int;
    reg PRLD_int;

//--------   JTAG Globals --------------
    wire JTAG_TDO_GLBL;
    wire JTAG_TCK_GLBL;
    wire JTAG_TDI_GLBL;
    wire JTAG_TMS_GLBL;
    wire JTAG_TRST_GLBL;

    reg JTAG_CAPTURE_GLBL;
    reg JTAG_RESET_GLBL;
    reg JTAG_SHIFT_GLBL;
    reg JTAG_UPDATE_GLBL;
    reg JTAG_RUNTEST_GLBL;

    reg JTAG_SEL1_GLBL = 0;
    reg JTAG_SEL2_GLBL = 0 ;
    reg JTAG_SEL3_GLBL = 0;
    reg JTAG_SEL4_GLBL = 0;

    reg JTAG_USER_TDO1_GLBL = 1'bz;
    reg JTAG_USER_TDO2_GLBL = 1'bz;
    reg JTAG_USER_TDO3_GLBL = 1'bz;
    reg JTAG_USER_TDO4_GLBL = 1'bz;

    assign (strong1, weak0) GSR = GSR_int;
    assign (strong1, weak0) GTS = GTS_int;
    assign (weak1, weak0) PRLD = PRLD_int;

    initial begin
	GSR_int = 1'b1;
	PRLD_int = 1'b1;
	#(ROC_WIDTH)
	GSR_int = 1'b0;
	PRLD_int = 1'b0;
    end

    initial begin
	GTS_int = 1'b1;
	#(TOC_WIDTH)
	GTS_int = 1'b0;
    end

endmodule
`endif
